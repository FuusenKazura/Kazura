module BranchPredictor(
  input         clock,
  input         reset,
  input  [15:0] io_pc,
  input         io_stall,
  input         io_learning_valid,
  input  [15:0] io_learning_bits_pc,
  input         io_learning_bits_result,
  output        io_predict
);
  reg [1:0] table_ [0:31]; // @[BranchPredictor.scala 27:35]
  reg [31:0] _RAND_0;
  wire [1:0] table___T_1_data; // @[BranchPredictor.scala 27:35]
  wire [4:0] table___T_1_addr; // @[BranchPredictor.scala 27:35]
  wire [1:0] table___T_25_data; // @[BranchPredictor.scala 27:35]
  wire [4:0] table___T_25_addr; // @[BranchPredictor.scala 27:35]
  wire [1:0] table___T_22_data; // @[BranchPredictor.scala 27:35]
  wire [4:0] table___T_22_addr; // @[BranchPredictor.scala 27:35]
  wire  table___T_22_mask; // @[BranchPredictor.scala 27:35]
  wire  table___T_22_en; // @[BranchPredictor.scala 27:35]
  reg [15:0] prev_pc; // @[BranchPredictor.scala 49:30]
  reg [31:0] _RAND_1;
  wire [15:0] pc; // @[BranchPredictor.scala 50:21]
  reg [15:0] addr; // @[BranchPredictor.scala 55:27]
  reg [31:0] _RAND_2;
  wire  _T_2; // @[Mux.scala 68:19]
  wire  _T_4; // @[Mux.scala 68:19]
  wire  _T_6; // @[Mux.scala 68:19]
  wire  _T_8; // @[Mux.scala 68:19]
  reg [1:0] updated; // @[BranchPredictor.scala 56:30]
  reg [31:0] _RAND_3;
  reg  _T_19; // @[BranchPredictor.scala 57:16]
  reg [31:0] _RAND_4;
  wire  _T_30; // @[Mux.scala 68:19]
  wire  _T_31; // @[Mux.scala 68:16]
  wire  _T_32; // @[Mux.scala 68:19]
  assign table___T_1_addr = io_learning_bits_pc[4:0];
  assign table___T_1_data = table_[table___T_1_addr]; // @[BranchPredictor.scala 27:35]
  assign table___T_25_addr = pc[4:0];
  assign table___T_25_data = table_[table___T_25_addr]; // @[BranchPredictor.scala 27:35]
  assign table___T_22_data = updated;
  assign table___T_22_addr = addr[4:0];
  assign table___T_22_mask = 1'h1;
  assign table___T_22_en = _T_19;
  assign pc = io_stall ? prev_pc : io_pc; // @[BranchPredictor.scala 50:21]
  assign _T_2 = 2'h3 == table___T_1_data; // @[Mux.scala 68:19]
  assign _T_4 = 2'h2 == table___T_1_data; // @[Mux.scala 68:19]
  assign _T_6 = 2'h1 == table___T_1_data; // @[Mux.scala 68:19]
  assign _T_8 = 2'h0 == table___T_1_data; // @[Mux.scala 68:19]
  assign _T_30 = 2'h1 == table___T_25_data; // @[Mux.scala 68:19]
  assign _T_31 = _T_30 ? 1'h0 : 1'h1; // @[Mux.scala 68:16]
  assign _T_32 = 2'h0 == table___T_25_data; // @[Mux.scala 68:19]
  assign io_predict = _T_32 ? 1'h0 : _T_31; // @[BranchPredictor.scala 61:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    table_[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  prev_pc = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  updated = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_19 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(table___T_22_en & table___T_22_mask) begin
      table_[table___T_22_addr] <= table___T_22_data; // @[BranchPredictor.scala 27:35]
    end
    if (reset) begin
      prev_pc <= io_pc;
    end else if (!(io_stall)) begin
      prev_pc <= io_pc;
    end
    addr <= io_learning_bits_pc;
    if (io_learning_bits_result) begin
      if (_T_8) begin
        updated <= 2'h1;
      end else if (_T_6) begin
        updated <= 2'h2;
      end else if (_T_4) begin
        updated <= 2'h3;
      end else if (_T_2) begin
        updated <= 2'h3;
      end else begin
        updated <= 2'h0;
      end
    end else if (_T_8) begin
      updated <= 2'h0;
    end else if (_T_6) begin
      updated <= 2'h0;
    end else if (_T_4) begin
      updated <= 2'h1;
    end else if (_T_2) begin
      updated <= 2'h2;
    end else begin
      updated <= 2'h0;
    end
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= io_learning_valid;
    end
  end
endmodule
module Fetch(
  input         clock,
  input         reset,
  input  [15:0] io_prev_pc,
  input         io_in_branch_mispredicted,
  input         io_in_branch_graduated,
  input  [15:0] io_in_restoration_pc,
  input         io_in_predict,
  input         io_in_predict_enable,
  input  [15:0] io_in_predict_pc,
  input         io_in_is_jump,
  input  [15:0] io_in_jump_pc,
  input         io_in_stall,
  output [15:0] io_out_pc
);
  wire [15:0] next_pc; // @[Fetch.scala 21:34]
  wire  _T_1; // @[Fetch.scala 25:29]
  wire  _T_2; // @[Fetch.scala 29:27]
  wire [15:0] _T_3; // @[Mux.scala 87:16]
  wire [15:0] _T_4; // @[Mux.scala 87:16]
  wire [15:0] _T_5; // @[Mux.scala 87:16]
  wire  _T_7; // @[Fetch.scala 34:9]
  wire  _T_8; // @[Fetch.scala 34:9]
  assign next_pc = io_prev_pc + 16'h1; // @[Fetch.scala 21:34]
  assign _T_1 = io_in_branch_graduated & io_in_branch_mispredicted; // @[Fetch.scala 25:29]
  assign _T_2 = io_in_predict_enable & io_in_predict; // @[Fetch.scala 29:27]
  assign _T_3 = io_in_stall ? io_prev_pc : next_pc; // @[Mux.scala 87:16]
  assign _T_4 = _T_2 ? io_in_predict_pc : _T_3; // @[Mux.scala 87:16]
  assign _T_5 = io_in_is_jump ? io_in_jump_pc : _T_4; // @[Mux.scala 87:16]
  assign _T_7 = $unsigned(reset); // @[Fetch.scala 34:9]
  assign _T_8 = _T_7 == 1'h0; // @[Fetch.scala 34:9]
  assign io_out_pc = _T_1 ? io_in_restoration_pc : _T_5; // @[Fetch.scala 23:13]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8) begin
          $fwrite(32'h80000002,"pc: %d, next_pc: %d, branch_mispredicted_enable: %d, branch_mispredicted: %d, restore_pc: %d\n",io_prev_pc,io_out_pc,io_in_branch_graduated,io_in_branch_mispredicted,io_in_restoration_pc); // @[Fetch.scala 34:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IF(
  input         clock,
  input         reset,
  input         io_in_branch_mispredicted,
  input         io_in_branch_graduated,
  input  [15:0] io_in_restoration_pc,
  input         io_in_predict,
  input         io_in_predict_enable,
  input  [15:0] io_in_predict_pc,
  input         io_in_is_jump,
  input  [15:0] io_in_jump_pc,
  input         io_in_stall,
  output [15:0] io_out_pc,
  output [15:0] io_out_total_cnt,
  output [3:0]  io_out_inst_bits_op,
  output [2:0]  io_out_inst_bits_rd,
  output [2:0]  io_out_inst_bits_rs,
  output [5:0]  io_out_inst_bits_disp6u
);
  wire  fetch_clock; // @[IF.scala 39:28]
  wire  fetch_reset; // @[IF.scala 39:28]
  wire [15:0] fetch_io_prev_pc; // @[IF.scala 39:28]
  wire  fetch_io_in_branch_mispredicted; // @[IF.scala 39:28]
  wire  fetch_io_in_branch_graduated; // @[IF.scala 39:28]
  wire [15:0] fetch_io_in_restoration_pc; // @[IF.scala 39:28]
  wire  fetch_io_in_predict; // @[IF.scala 39:28]
  wire  fetch_io_in_predict_enable; // @[IF.scala 39:28]
  wire [15:0] fetch_io_in_predict_pc; // @[IF.scala 39:28]
  wire  fetch_io_in_is_jump; // @[IF.scala 39:28]
  wire [15:0] fetch_io_in_jump_pc; // @[IF.scala 39:28]
  wire  fetch_io_in_stall; // @[IF.scala 39:28]
  wire [15:0] fetch_io_out_pc; // @[IF.scala 39:28]
  reg [15:0] pc; // @[IF.scala 35:25]
  reg [31:0] _RAND_0;
  reg [15:0] total_cnt; // @[IF.scala 36:32]
  reg [31:0] _RAND_1;
  wire [15:0] _T_2; // @[IF.scala 37:26]
  wire [4:0] _T_3;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_4;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  Fetch fetch ( // @[IF.scala 39:28]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_prev_pc(fetch_io_prev_pc),
    .io_in_branch_mispredicted(fetch_io_in_branch_mispredicted),
    .io_in_branch_graduated(fetch_io_in_branch_graduated),
    .io_in_restoration_pc(fetch_io_in_restoration_pc),
    .io_in_predict(fetch_io_in_predict),
    .io_in_predict_enable(fetch_io_in_predict_enable),
    .io_in_predict_pc(fetch_io_in_predict_pc),
    .io_in_is_jump(fetch_io_in_is_jump),
    .io_in_jump_pc(fetch_io_in_jump_pc),
    .io_in_stall(fetch_io_in_stall),
    .io_out_pc(fetch_io_out_pc)
  );
  assign _T_2 = total_cnt + 16'h1; // @[IF.scala 37:26]
  assign _T_3 = pc[4:0];
  assign _GEN_1 = 5'h1 == _T_3 ? 16'h9400 : 16'h9200;
  assign _GEN_2 = 5'h2 == _T_3 ? 16'h9609 : _GEN_1;
  assign _GEN_3 = 5'h3 == _T_3 ? 16'h9800 : _GEN_2;
  assign _GEN_4 = 5'h4 == _T_3 ? 16'h5201 : _GEN_3;
  assign _GEN_5 = 5'h5 == _T_3 ? 16'h1440 : _GEN_4;
  assign _GEN_6 = 5'h6 == _T_3 ? 16'hd2c3 : _GEN_5;
  assign _GEN_7 = 5'h7 == _T_3 ? 16'h0 : _GEN_6;
  assign _GEN_8 = 5'h8 == _T_3 ? 16'he1fc : _GEN_7;
  assign _GEN_9 = 5'h9 == _T_3 ? 16'h1880 : _GEN_8;
  assign _GEN_10 = 5'ha == _T_3 ? 16'h0 : _GEN_9;
  assign _GEN_11 = 5'hb == _T_3 ? 16'h0 : _GEN_10;
  assign _GEN_12 = 5'hc == _T_3 ? 16'h0 : _GEN_11;
  assign _GEN_13 = 5'hd == _T_3 ? 16'h0 : _GEN_12;
  assign _GEN_14 = 5'he == _T_3 ? 16'h0 : _GEN_13;
  assign _GEN_15 = 5'hf == _T_3 ? 16'h0 : _GEN_14;
  assign _GEN_16 = 5'h10 == _T_3 ? 16'h0 : _GEN_15;
  assign _GEN_17 = 5'h11 == _T_3 ? 16'h0 : _GEN_16;
  assign _GEN_18 = 5'h12 == _T_3 ? 16'h0 : _GEN_17;
  assign _GEN_19 = 5'h13 == _T_3 ? 16'h0 : _GEN_18;
  assign _GEN_20 = 5'h14 == _T_3 ? 16'h0 : _GEN_19;
  assign _GEN_21 = 5'h15 == _T_3 ? 16'h0 : _GEN_20;
  assign _GEN_22 = 5'h16 == _T_3 ? 16'h0 : _GEN_21;
  assign _GEN_23 = 5'h17 == _T_3 ? 16'h0 : _GEN_22;
  assign _GEN_24 = 5'h18 == _T_3 ? 16'h0 : _GEN_23;
  assign _GEN_25 = 5'h19 == _T_3 ? 16'h0 : _GEN_24;
  assign _GEN_26 = 5'h1a == _T_3 ? 16'h0 : _GEN_25;
  assign _GEN_27 = 5'h1b == _T_3 ? 16'h0 : _GEN_26;
  assign _GEN_28 = 5'h1c == _T_3 ? 16'h0 : _GEN_27;
  assign _GEN_29 = 5'h1d == _T_3 ? 16'h0 : _GEN_28;
  assign _GEN_30 = 5'h1e == _T_3 ? 16'h0 : _GEN_29;
  assign _GEN_31 = 5'h1f == _T_3 ? 16'h0 : _GEN_30;
  assign io_out_pc = pc; // @[IF.scala 55:13]
  assign io_out_total_cnt = total_cnt; // @[IF.scala 56:20]
  assign io_out_inst_bits_op = _GEN_31[15:12]; // @[IF.scala 57:20]
  assign io_out_inst_bits_rd = _GEN_31[11:9]; // @[IF.scala 57:20]
  assign io_out_inst_bits_rs = _GEN_31[8:6]; // @[IF.scala 57:20]
  assign io_out_inst_bits_disp6u = _GEN_31[5:0]; // @[IF.scala 57:20]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_prev_pc = pc; // @[IF.scala 51:20]
  assign fetch_io_in_branch_mispredicted = io_in_branch_mispredicted; // @[IF.scala 43:35]
  assign fetch_io_in_branch_graduated = io_in_branch_graduated; // @[IF.scala 44:32]
  assign fetch_io_in_restoration_pc = io_in_restoration_pc; // @[IF.scala 45:30]
  assign fetch_io_in_predict = io_in_predict; // @[IF.scala 40:23]
  assign fetch_io_in_predict_enable = io_in_predict_enable; // @[IF.scala 41:30]
  assign fetch_io_in_predict_pc = io_in_predict_pc; // @[IF.scala 42:26]
  assign fetch_io_in_is_jump = io_in_is_jump; // @[IF.scala 47:23]
  assign fetch_io_in_jump_pc = io_in_jump_pc; // @[IF.scala 48:23]
  assign fetch_io_in_stall = io_in_stall; // @[IF.scala 49:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  total_cnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 16'h0;
    end else begin
      pc <= fetch_io_out_pc;
    end
    if (reset) begin
      total_cnt <= 16'h0;
    end else begin
      total_cnt <= _T_2;
    end
  end
endmodule
module Decoder(
  input  [3:0]  io_inst_bits_op,
  output [2:0]  io_ctrl_alu_op,
  output        io_ctrl_is_jump,
  output        io_ctrl_is_branch,
  output        io_ctrl_rf_w,
  output        io_ctrl_mem_r,
  output        io_ctrl_mem_w,
  output        io_ctrl_rs1_use,
  output        io_ctrl_rs2_use,
  output [15:0] io_source_sel_0,
  output [15:0] io_source_sel_1
);
  wire  _T; // @[Decoder.scala 36:26]
  wire  _T_1; // @[Decoder.scala 39:32]
  wire  _T_2; // @[Decoder.scala 39:32]
  wire  _T_3; // @[Decoder.scala 39:32]
  wire  _T_4; // @[Decoder.scala 39:32]
  wire  _T_5; // @[Decoder.scala 39:32]
  wire  _T_6; // @[Decoder.scala 39:32]
  wire  _T_7; // @[Decoder.scala 39:32]
  wire  _T_9; // @[Decoder.scala 39:32]
  wire  _T_10; // @[Decoder.scala 39:32]
  wire  _T_11; // @[Decoder.scala 39:32]
  wire  _T_12; // @[Decoder.scala 39:32]
  wire  _T_13; // @[Decoder.scala 39:32]
  wire  _T_14; // @[Decoder.scala 39:32]
  wire  _T_15; // @[Decoder.scala 39:32]
  wire [1:0] _GEN_3; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_4; // @[Decoder.scala 39:45]
  wire  _GEN_5; // @[Decoder.scala 39:45]
  wire  _GEN_8; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_9; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_10; // @[Decoder.scala 39:45]
  wire  _GEN_11; // @[Decoder.scala 39:45]
  wire  _GEN_12; // @[Decoder.scala 39:45]
  wire  _GEN_14; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_15; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_16; // @[Decoder.scala 39:45]
  wire  _GEN_17; // @[Decoder.scala 39:45]
  wire  _GEN_18; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_21; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_22; // @[Decoder.scala 39:45]
  wire  _GEN_23; // @[Decoder.scala 39:45]
  wire  _GEN_24; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_25; // @[Decoder.scala 39:45]
  wire  _GEN_26; // @[Decoder.scala 39:45]
  wire  _GEN_27; // @[Decoder.scala 39:45]
  wire  _GEN_30; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_31; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_32; // @[Decoder.scala 39:45]
  wire  _GEN_33; // @[Decoder.scala 39:45]
  wire  _GEN_34; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_35; // @[Decoder.scala 39:45]
  wire  _GEN_36; // @[Decoder.scala 39:45]
  wire  _GEN_37; // @[Decoder.scala 39:45]
  wire  _GEN_39; // @[Decoder.scala 39:45]
  wire  _GEN_40; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_41; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_42; // @[Decoder.scala 39:45]
  wire  _GEN_43; // @[Decoder.scala 39:45]
  wire  _GEN_44; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_45; // @[Decoder.scala 39:45]
  wire  _GEN_46; // @[Decoder.scala 39:45]
  wire  _GEN_47; // @[Decoder.scala 39:45]
  wire  _GEN_48; // @[Decoder.scala 39:45]
  wire  _GEN_49; // @[Decoder.scala 39:45]
  wire  _GEN_50; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_51; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_52; // @[Decoder.scala 39:45]
  wire  _GEN_53; // @[Decoder.scala 39:45]
  wire  _GEN_54; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_55; // @[Decoder.scala 39:45]
  wire  _GEN_56; // @[Decoder.scala 39:45]
  wire  _GEN_57; // @[Decoder.scala 39:45]
  wire  _GEN_58; // @[Decoder.scala 39:45]
  wire  _GEN_59; // @[Decoder.scala 39:45]
  wire  _GEN_60; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_61; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_62; // @[Decoder.scala 39:45]
  wire  _GEN_63; // @[Decoder.scala 39:45]
  wire  _GEN_64; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_65; // @[Decoder.scala 39:45]
  wire  _GEN_66; // @[Decoder.scala 39:45]
  wire  _GEN_67; // @[Decoder.scala 39:45]
  wire  _GEN_68; // @[Decoder.scala 39:45]
  wire  _GEN_69; // @[Decoder.scala 39:45]
  wire  _GEN_70; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_71; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_72; // @[Decoder.scala 39:45]
  wire  _GEN_73; // @[Decoder.scala 39:45]
  wire  _GEN_74; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_75; // @[Decoder.scala 39:45]
  wire  _GEN_76; // @[Decoder.scala 39:45]
  wire  _GEN_77; // @[Decoder.scala 39:45]
  wire  _GEN_78; // @[Decoder.scala 39:45]
  wire  _GEN_79; // @[Decoder.scala 39:45]
  wire  _GEN_80; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_81; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_82; // @[Decoder.scala 39:45]
  wire  _GEN_83; // @[Decoder.scala 39:45]
  wire  _GEN_84; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_85; // @[Decoder.scala 39:45]
  wire  _GEN_86; // @[Decoder.scala 39:45]
  wire  _GEN_87; // @[Decoder.scala 39:45]
  wire  _GEN_88; // @[Decoder.scala 39:45]
  wire  _GEN_89; // @[Decoder.scala 39:45]
  wire  _GEN_90; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_91; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_92; // @[Decoder.scala 39:45]
  wire  _GEN_93; // @[Decoder.scala 39:45]
  wire  _GEN_94; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_95; // @[Decoder.scala 39:45]
  wire  _GEN_96; // @[Decoder.scala 39:45]
  wire  _GEN_97; // @[Decoder.scala 39:45]
  wire  _GEN_98; // @[Decoder.scala 39:45]
  wire  _GEN_99; // @[Decoder.scala 39:45]
  wire  _GEN_100; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_101; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_102; // @[Decoder.scala 39:45]
  wire  _GEN_103; // @[Decoder.scala 39:45]
  wire  _GEN_104; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_105; // @[Decoder.scala 39:45]
  wire  _GEN_106; // @[Decoder.scala 39:45]
  wire  _GEN_107; // @[Decoder.scala 39:45]
  wire  _GEN_108; // @[Decoder.scala 39:45]
  wire  _GEN_109; // @[Decoder.scala 39:45]
  wire  _GEN_110; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_111; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_112; // @[Decoder.scala 39:45]
  wire  _GEN_113; // @[Decoder.scala 39:45]
  wire  _GEN_114; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_115; // @[Decoder.scala 39:45]
  wire  _GEN_116; // @[Decoder.scala 39:45]
  wire  _GEN_117; // @[Decoder.scala 39:45]
  wire  _GEN_118; // @[Decoder.scala 39:45]
  wire  _GEN_119; // @[Decoder.scala 39:45]
  wire  _GEN_120; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_121; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_122; // @[Decoder.scala 39:45]
  wire  _GEN_123; // @[Decoder.scala 39:45]
  wire  _GEN_124; // @[Decoder.scala 39:45]
  wire [2:0] _GEN_125; // @[Decoder.scala 39:45]
  wire  _GEN_126; // @[Decoder.scala 39:45]
  wire  _GEN_127; // @[Decoder.scala 39:45]
  wire  _GEN_128; // @[Decoder.scala 39:45]
  wire  _GEN_129; // @[Decoder.scala 39:45]
  wire  _GEN_130; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_131; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_132; // @[Decoder.scala 39:45]
  wire  _GEN_133; // @[Decoder.scala 39:45]
  wire  _GEN_134; // @[Decoder.scala 39:45]
  wire [1:0] _GEN_141; // @[Decoder.scala 36:38]
  wire [1:0] _GEN_142; // @[Decoder.scala 36:38]
  assign _T = io_inst_bits_op == 4'h0; // @[Decoder.scala 36:26]
  assign _T_1 = io_inst_bits_op == 4'h1; // @[Decoder.scala 39:32]
  assign _T_2 = io_inst_bits_op == 4'h2; // @[Decoder.scala 39:32]
  assign _T_3 = io_inst_bits_op == 4'h3; // @[Decoder.scala 39:32]
  assign _T_4 = io_inst_bits_op == 4'h4; // @[Decoder.scala 39:32]
  assign _T_5 = io_inst_bits_op == 4'h5; // @[Decoder.scala 39:32]
  assign _T_6 = io_inst_bits_op == 4'h6; // @[Decoder.scala 39:32]
  assign _T_7 = io_inst_bits_op == 4'h7; // @[Decoder.scala 39:32]
  assign _T_9 = io_inst_bits_op == 4'h8; // @[Decoder.scala 39:32]
  assign _T_10 = io_inst_bits_op == 4'h9; // @[Decoder.scala 39:32]
  assign _T_11 = io_inst_bits_op == 4'ha; // @[Decoder.scala 39:32]
  assign _T_12 = io_inst_bits_op == 4'hb; // @[Decoder.scala 39:32]
  assign _T_13 = io_inst_bits_op == 4'hc; // @[Decoder.scala 39:32]
  assign _T_14 = io_inst_bits_op == 4'hd; // @[Decoder.scala 39:32]
  assign _T_15 = io_inst_bits_op == 4'he; // @[Decoder.scala 39:32]
  assign _GEN_3 = _T_15 ? 2'h2 : 2'h0; // @[Decoder.scala 39:45]
  assign _GEN_4 = _T_14 ? 3'h5 : 3'h0; // @[Decoder.scala 39:45]
  assign _GEN_5 = _T_14 ? 1'h0 : _T_15; // @[Decoder.scala 39:45]
  assign _GEN_8 = _T_14 | _T_15; // @[Decoder.scala 39:45]
  assign _GEN_9 = _T_14 ? 2'h1 : _GEN_3; // @[Decoder.scala 39:45]
  assign _GEN_10 = _T_13 ? 3'h4 : _GEN_4; // @[Decoder.scala 39:45]
  assign _GEN_11 = _T_13 ? 1'h0 : _GEN_5; // @[Decoder.scala 39:45]
  assign _GEN_12 = _T_13 | _T_14; // @[Decoder.scala 39:45]
  assign _GEN_14 = _T_13 | _GEN_8; // @[Decoder.scala 39:45]
  assign _GEN_15 = _T_13 ? 2'h1 : _GEN_9; // @[Decoder.scala 39:45]
  assign _GEN_16 = _T_12 ? 3'h0 : _GEN_10; // @[Decoder.scala 39:45]
  assign _GEN_17 = _T_12 ? 1'h0 : _GEN_11; // @[Decoder.scala 39:45]
  assign _GEN_18 = _T_12 ? 1'h0 : _GEN_12; // @[Decoder.scala 39:45]
  assign _GEN_21 = _T_12 ? 2'h3 : {{1'd0}, _GEN_14}; // @[Decoder.scala 39:45]
  assign _GEN_22 = _T_12 ? 2'h1 : _GEN_15; // @[Decoder.scala 39:45]
  assign _GEN_23 = _T_12 | _GEN_14; // @[Decoder.scala 39:45]
  assign _GEN_24 = _T_12 | _GEN_12; // @[Decoder.scala 39:45]
  assign _GEN_25 = _T_11 ? 3'h0 : _GEN_16; // @[Decoder.scala 39:45]
  assign _GEN_26 = _T_11 ? 1'h0 : _GEN_17; // @[Decoder.scala 39:45]
  assign _GEN_27 = _T_11 ? 1'h0 : _GEN_18; // @[Decoder.scala 39:45]
  assign _GEN_30 = _T_11 ? 1'h0 : _T_12; // @[Decoder.scala 39:45]
  assign _GEN_31 = _T_11 ? 2'h3 : _GEN_21; // @[Decoder.scala 39:45]
  assign _GEN_32 = _T_11 ? 2'h1 : _GEN_22; // @[Decoder.scala 39:45]
  assign _GEN_33 = _T_11 ? 1'h0 : _GEN_23; // @[Decoder.scala 39:45]
  assign _GEN_34 = _T_11 | _GEN_24; // @[Decoder.scala 39:45]
  assign _GEN_35 = _T_10 ? 3'h0 : _GEN_25; // @[Decoder.scala 39:45]
  assign _GEN_36 = _T_10 ? 1'h0 : _GEN_26; // @[Decoder.scala 39:45]
  assign _GEN_37 = _T_10 ? 1'h0 : _GEN_27; // @[Decoder.scala 39:45]
  assign _GEN_39 = _T_10 ? 1'h0 : _T_11; // @[Decoder.scala 39:45]
  assign _GEN_40 = _T_10 ? 1'h0 : _GEN_30; // @[Decoder.scala 39:45]
  assign _GEN_41 = _T_10 ? 2'h0 : _GEN_31; // @[Decoder.scala 39:45]
  assign _GEN_42 = _T_10 ? 2'h2 : _GEN_32; // @[Decoder.scala 39:45]
  assign _GEN_43 = _T_10 ? 1'h0 : _GEN_33; // @[Decoder.scala 39:45]
  assign _GEN_44 = _T_10 ? 1'h0 : _GEN_34; // @[Decoder.scala 39:45]
  assign _GEN_45 = _T_9 ? 3'h1 : _GEN_35; // @[Decoder.scala 39:45]
  assign _GEN_46 = _T_9 ? 1'h0 : _GEN_36; // @[Decoder.scala 39:45]
  assign _GEN_47 = _T_9 ? 1'h0 : _GEN_37; // @[Decoder.scala 39:45]
  assign _GEN_48 = _T_9 | _T_10; // @[Decoder.scala 39:45]
  assign _GEN_49 = _T_9 ? 1'h0 : _GEN_39; // @[Decoder.scala 39:45]
  assign _GEN_50 = _T_9 ? 1'h0 : _GEN_40; // @[Decoder.scala 39:45]
  assign _GEN_51 = _T_9 ? 2'h1 : _GEN_41; // @[Decoder.scala 39:45]
  assign _GEN_52 = _T_9 ? 2'h0 : _GEN_42; // @[Decoder.scala 39:45]
  assign _GEN_53 = _T_9 | _GEN_43; // @[Decoder.scala 39:45]
  assign _GEN_54 = _T_9 ? 1'h0 : _GEN_44; // @[Decoder.scala 39:45]
  assign _GEN_55 = _T_7 ? 3'h0 : _GEN_45; // @[Decoder.scala 39:45]
  assign _GEN_56 = _T_7 ? 1'h0 : _GEN_46; // @[Decoder.scala 39:45]
  assign _GEN_57 = _T_7 ? 1'h0 : _GEN_47; // @[Decoder.scala 39:45]
  assign _GEN_58 = _T_7 | _GEN_48; // @[Decoder.scala 39:45]
  assign _GEN_59 = _T_7 ? 1'h0 : _GEN_49; // @[Decoder.scala 39:45]
  assign _GEN_60 = _T_7 ? 1'h0 : _GEN_50; // @[Decoder.scala 39:45]
  assign _GEN_61 = _T_7 ? 2'h1 : _GEN_51; // @[Decoder.scala 39:45]
  assign _GEN_62 = _T_7 ? 2'h0 : _GEN_52; // @[Decoder.scala 39:45]
  assign _GEN_63 = _T_7 | _GEN_53; // @[Decoder.scala 39:45]
  assign _GEN_64 = _T_7 ? 1'h0 : _GEN_54; // @[Decoder.scala 39:45]
  assign _GEN_65 = _T_7 ? 3'h0 : _GEN_55; // @[Decoder.scala 39:45]
  assign _GEN_66 = _T_7 ? 1'h0 : _GEN_56; // @[Decoder.scala 39:45]
  assign _GEN_67 = _T_7 ? 1'h0 : _GEN_57; // @[Decoder.scala 39:45]
  assign _GEN_68 = _T_7 | _GEN_58; // @[Decoder.scala 39:45]
  assign _GEN_69 = _T_7 ? 1'h0 : _GEN_59; // @[Decoder.scala 39:45]
  assign _GEN_70 = _T_7 ? 1'h0 : _GEN_60; // @[Decoder.scala 39:45]
  assign _GEN_71 = _T_7 ? 2'h1 : _GEN_61; // @[Decoder.scala 39:45]
  assign _GEN_72 = _T_7 ? 2'h0 : _GEN_62; // @[Decoder.scala 39:45]
  assign _GEN_73 = _T_7 | _GEN_63; // @[Decoder.scala 39:45]
  assign _GEN_74 = _T_7 ? 1'h0 : _GEN_64; // @[Decoder.scala 39:45]
  assign _GEN_75 = _T_6 ? 3'h1 : _GEN_65; // @[Decoder.scala 39:45]
  assign _GEN_76 = _T_6 ? 1'h0 : _GEN_66; // @[Decoder.scala 39:45]
  assign _GEN_77 = _T_6 ? 1'h0 : _GEN_67; // @[Decoder.scala 39:45]
  assign _GEN_78 = _T_6 | _GEN_68; // @[Decoder.scala 39:45]
  assign _GEN_79 = _T_6 ? 1'h0 : _GEN_69; // @[Decoder.scala 39:45]
  assign _GEN_80 = _T_6 ? 1'h0 : _GEN_70; // @[Decoder.scala 39:45]
  assign _GEN_81 = _T_6 ? 2'h1 : _GEN_71; // @[Decoder.scala 39:45]
  assign _GEN_82 = _T_6 ? 2'h2 : _GEN_72; // @[Decoder.scala 39:45]
  assign _GEN_83 = _T_6 | _GEN_73; // @[Decoder.scala 39:45]
  assign _GEN_84 = _T_6 ? 1'h0 : _GEN_74; // @[Decoder.scala 39:45]
  assign _GEN_85 = _T_5 ? 3'h0 : _GEN_75; // @[Decoder.scala 39:45]
  assign _GEN_86 = _T_5 ? 1'h0 : _GEN_76; // @[Decoder.scala 39:45]
  assign _GEN_87 = _T_5 ? 1'h0 : _GEN_77; // @[Decoder.scala 39:45]
  assign _GEN_88 = _T_5 | _GEN_78; // @[Decoder.scala 39:45]
  assign _GEN_89 = _T_5 ? 1'h0 : _GEN_79; // @[Decoder.scala 39:45]
  assign _GEN_90 = _T_5 ? 1'h0 : _GEN_80; // @[Decoder.scala 39:45]
  assign _GEN_91 = _T_5 ? 2'h1 : _GEN_81; // @[Decoder.scala 39:45]
  assign _GEN_92 = _T_5 ? 2'h2 : _GEN_82; // @[Decoder.scala 39:45]
  assign _GEN_93 = _T_5 | _GEN_83; // @[Decoder.scala 39:45]
  assign _GEN_94 = _T_5 ? 1'h0 : _GEN_84; // @[Decoder.scala 39:45]
  assign _GEN_95 = _T_4 ? 3'h3 : _GEN_85; // @[Decoder.scala 39:45]
  assign _GEN_96 = _T_4 ? 1'h0 : _GEN_86; // @[Decoder.scala 39:45]
  assign _GEN_97 = _T_4 ? 1'h0 : _GEN_87; // @[Decoder.scala 39:45]
  assign _GEN_98 = _T_4 | _GEN_88; // @[Decoder.scala 39:45]
  assign _GEN_99 = _T_4 ? 1'h0 : _GEN_89; // @[Decoder.scala 39:45]
  assign _GEN_100 = _T_4 ? 1'h0 : _GEN_90; // @[Decoder.scala 39:45]
  assign _GEN_101 = _T_4 ? 2'h1 : _GEN_91; // @[Decoder.scala 39:45]
  assign _GEN_102 = _T_4 ? 2'h1 : _GEN_92; // @[Decoder.scala 39:45]
  assign _GEN_103 = _T_4 | _GEN_93; // @[Decoder.scala 39:45]
  assign _GEN_104 = _T_4 | _GEN_94; // @[Decoder.scala 39:45]
  assign _GEN_105 = _T_3 ? 3'h2 : _GEN_95; // @[Decoder.scala 39:45]
  assign _GEN_106 = _T_3 ? 1'h0 : _GEN_96; // @[Decoder.scala 39:45]
  assign _GEN_107 = _T_3 ? 1'h0 : _GEN_97; // @[Decoder.scala 39:45]
  assign _GEN_108 = _T_3 | _GEN_98; // @[Decoder.scala 39:45]
  assign _GEN_109 = _T_3 ? 1'h0 : _GEN_99; // @[Decoder.scala 39:45]
  assign _GEN_110 = _T_3 ? 1'h0 : _GEN_100; // @[Decoder.scala 39:45]
  assign _GEN_111 = _T_3 ? 2'h1 : _GEN_101; // @[Decoder.scala 39:45]
  assign _GEN_112 = _T_3 ? 2'h1 : _GEN_102; // @[Decoder.scala 39:45]
  assign _GEN_113 = _T_3 | _GEN_103; // @[Decoder.scala 39:45]
  assign _GEN_114 = _T_3 | _GEN_104; // @[Decoder.scala 39:45]
  assign _GEN_115 = _T_2 ? 3'h1 : _GEN_105; // @[Decoder.scala 39:45]
  assign _GEN_116 = _T_2 ? 1'h0 : _GEN_106; // @[Decoder.scala 39:45]
  assign _GEN_117 = _T_2 ? 1'h0 : _GEN_107; // @[Decoder.scala 39:45]
  assign _GEN_118 = _T_2 | _GEN_108; // @[Decoder.scala 39:45]
  assign _GEN_119 = _T_2 ? 1'h0 : _GEN_109; // @[Decoder.scala 39:45]
  assign _GEN_120 = _T_2 ? 1'h0 : _GEN_110; // @[Decoder.scala 39:45]
  assign _GEN_121 = _T_2 ? 2'h1 : _GEN_111; // @[Decoder.scala 39:45]
  assign _GEN_122 = _T_2 ? 2'h1 : _GEN_112; // @[Decoder.scala 39:45]
  assign _GEN_123 = _T_2 | _GEN_113; // @[Decoder.scala 39:45]
  assign _GEN_124 = _T_2 | _GEN_114; // @[Decoder.scala 39:45]
  assign _GEN_125 = _T_1 ? 3'h0 : _GEN_115; // @[Decoder.scala 39:45]
  assign _GEN_126 = _T_1 ? 1'h0 : _GEN_116; // @[Decoder.scala 39:45]
  assign _GEN_127 = _T_1 ? 1'h0 : _GEN_117; // @[Decoder.scala 39:45]
  assign _GEN_128 = _T_1 | _GEN_118; // @[Decoder.scala 39:45]
  assign _GEN_129 = _T_1 ? 1'h0 : _GEN_119; // @[Decoder.scala 39:45]
  assign _GEN_130 = _T_1 ? 1'h0 : _GEN_120; // @[Decoder.scala 39:45]
  assign _GEN_131 = _T_1 ? 2'h1 : _GEN_121; // @[Decoder.scala 39:45]
  assign _GEN_132 = _T_1 ? 2'h1 : _GEN_122; // @[Decoder.scala 39:45]
  assign _GEN_133 = _T_1 | _GEN_123; // @[Decoder.scala 39:45]
  assign _GEN_134 = _T_1 | _GEN_124; // @[Decoder.scala 39:45]
  assign _GEN_141 = _T ? 2'h0 : _GEN_131; // @[Decoder.scala 36:38]
  assign _GEN_142 = _T ? 2'h0 : _GEN_132; // @[Decoder.scala 36:38]
  assign io_ctrl_alu_op = _T ? 3'h0 : _GEN_125; // @[Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23 Decoder.scala 21:23]
  assign io_ctrl_is_jump = _T ? 1'h0 : _GEN_126; // @[Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23 Decoder.scala 22:23]
  assign io_ctrl_is_branch = _T ? 1'h0 : _GEN_127; // @[Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23 Decoder.scala 23:23]
  assign io_ctrl_rf_w = _T ? 1'h0 : _GEN_128; // @[Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23 Decoder.scala 24:23]
  assign io_ctrl_mem_r = _T ? 1'h0 : _GEN_129; // @[Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23 Decoder.scala 25:23]
  assign io_ctrl_mem_w = _T ? 1'h0 : _GEN_130; // @[Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23 Decoder.scala 26:23]
  assign io_ctrl_rs1_use = _T ? 1'h0 : _GEN_133; // @[Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24 Decoder.scala 30:24]
  assign io_ctrl_rs2_use = _T ? 1'h0 : _GEN_134; // @[Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24 Decoder.scala 31:24]
  assign io_source_sel_0 = {{14'd0}, _GEN_141}; // @[Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24]
  assign io_source_sel_1 = {{14'd0}, _GEN_142}; // @[Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24 Decoder.scala 28:24]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [2:0]  io_read_addr_0,
  input  [2:0]  io_read_addr_1,
  input  [2:0]  io_write_0_rd_addr,
  input         io_write_0_rf_w,
  input  [15:0] io_write_0_data,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_rf4debug_1,
  output [15:0] io_rf4debug_2,
  output [15:0] io_rf4debug_3,
  output [15:0] io_rf4debug_4,
  output [15:0] io_rf4debug_5,
  output [15:0] io_rf4debug_6,
  output [15:0] io_rf4debug_7
);
  reg [15:0] rf_1; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_0;
  reg [15:0] rf_2; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_1;
  reg [15:0] rf_3; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_2;
  reg [15:0] rf_4; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_3;
  reg [15:0] rf_5; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_4;
  reg [15:0] rf_6; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_5;
  reg [15:0] rf_7; // @[RegisterFile.scala 23:26]
  reg [31:0] _RAND_6;
  wire  _T; // @[RegisterFile.scala 32:33]
  wire  _T_1; // @[RegisterFile.scala 32:19]
  wire [2:0] _T_2_rd_addr; // @[RegisterFile.scala 32:10]
  wire  _T_2_rf_w; // @[RegisterFile.scala 32:10]
  wire [15:0] _T_2_data; // @[RegisterFile.scala 32:10]
  wire  _T_4; // @[RegisterFile.scala 33:65]
  wire  _T_5; // @[RegisterFile.scala 33:40]
  wire [15:0] _GEN_1; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_2; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_3; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_4; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_5; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_6; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_7; // @[RegisterFile.scala 33:21]
  wire  _T_7; // @[RegisterFile.scala 32:33]
  wire  _T_8; // @[RegisterFile.scala 32:19]
  wire [2:0] _T_9_rd_addr; // @[RegisterFile.scala 32:10]
  wire  _T_9_rf_w; // @[RegisterFile.scala 32:10]
  wire [15:0] _T_9_data; // @[RegisterFile.scala 32:10]
  wire  _T_11; // @[RegisterFile.scala 33:65]
  wire  _T_12; // @[RegisterFile.scala 33:40]
  wire [15:0] _GEN_9; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_10; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_11; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_12; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_13; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_14; // @[RegisterFile.scala 33:21]
  wire [15:0] _GEN_15; // @[RegisterFile.scala 33:21]
  wire  _T_14; // @[RegisterFile.scala 49:11]
  wire  _T_15; // @[RegisterFile.scala 49:11]
  assign _T = io_write_0_rd_addr == io_read_addr_0; // @[RegisterFile.scala 32:33]
  assign _T_1 = io_write_0_rf_w & _T; // @[RegisterFile.scala 32:19]
  assign _T_2_rd_addr = _T_1 ? io_write_0_rd_addr : 3'h0; // @[RegisterFile.scala 32:10]
  assign _T_2_rf_w = _T_1 & io_write_0_rf_w; // @[RegisterFile.scala 32:10]
  assign _T_2_data = _T_1 ? io_write_0_data : 16'h0; // @[RegisterFile.scala 32:10]
  assign _T_4 = _T_2_rd_addr == io_read_addr_0; // @[RegisterFile.scala 33:65]
  assign _T_5 = _T_2_rf_w & _T_4; // @[RegisterFile.scala 33:40]
  assign _GEN_1 = 3'h1 == io_read_addr_0 ? rf_1 : 16'h0; // @[RegisterFile.scala 33:21]
  assign _GEN_2 = 3'h2 == io_read_addr_0 ? rf_2 : _GEN_1; // @[RegisterFile.scala 33:21]
  assign _GEN_3 = 3'h3 == io_read_addr_0 ? rf_3 : _GEN_2; // @[RegisterFile.scala 33:21]
  assign _GEN_4 = 3'h4 == io_read_addr_0 ? rf_4 : _GEN_3; // @[RegisterFile.scala 33:21]
  assign _GEN_5 = 3'h5 == io_read_addr_0 ? rf_5 : _GEN_4; // @[RegisterFile.scala 33:21]
  assign _GEN_6 = 3'h6 == io_read_addr_0 ? rf_6 : _GEN_5; // @[RegisterFile.scala 33:21]
  assign _GEN_7 = 3'h7 == io_read_addr_0 ? rf_7 : _GEN_6; // @[RegisterFile.scala 33:21]
  assign _T_7 = io_write_0_rd_addr == io_read_addr_1; // @[RegisterFile.scala 32:33]
  assign _T_8 = io_write_0_rf_w & _T_7; // @[RegisterFile.scala 32:19]
  assign _T_9_rd_addr = _T_8 ? io_write_0_rd_addr : 3'h0; // @[RegisterFile.scala 32:10]
  assign _T_9_rf_w = _T_8 & io_write_0_rf_w; // @[RegisterFile.scala 32:10]
  assign _T_9_data = _T_8 ? io_write_0_data : 16'h0; // @[RegisterFile.scala 32:10]
  assign _T_11 = _T_9_rd_addr == io_read_addr_1; // @[RegisterFile.scala 33:65]
  assign _T_12 = _T_9_rf_w & _T_11; // @[RegisterFile.scala 33:40]
  assign _GEN_9 = 3'h1 == io_read_addr_1 ? rf_1 : 16'h0; // @[RegisterFile.scala 33:21]
  assign _GEN_10 = 3'h2 == io_read_addr_1 ? rf_2 : _GEN_9; // @[RegisterFile.scala 33:21]
  assign _GEN_11 = 3'h3 == io_read_addr_1 ? rf_3 : _GEN_10; // @[RegisterFile.scala 33:21]
  assign _GEN_12 = 3'h4 == io_read_addr_1 ? rf_4 : _GEN_11; // @[RegisterFile.scala 33:21]
  assign _GEN_13 = 3'h5 == io_read_addr_1 ? rf_5 : _GEN_12; // @[RegisterFile.scala 33:21]
  assign _GEN_14 = 3'h6 == io_read_addr_1 ? rf_6 : _GEN_13; // @[RegisterFile.scala 33:21]
  assign _GEN_15 = 3'h7 == io_read_addr_1 ? rf_7 : _GEN_14; // @[RegisterFile.scala 33:21]
  assign _T_14 = $unsigned(reset); // @[RegisterFile.scala 49:11]
  assign _T_15 = _T_14 == 1'h0; // @[RegisterFile.scala 49:11]
  assign io_out_0 = _T_5 ? _T_2_data : _GEN_7; // @[RegisterFile.scala 33:15]
  assign io_out_1 = _T_12 ? _T_9_data : _GEN_15; // @[RegisterFile.scala 33:15]
  assign io_rf4debug_1 = rf_1; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_2 = rf_2; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_3 = rf_3; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_4 = rf_4; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_5 = rf_5; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_6 = rf_6; // @[RegisterFile.scala 46:15]
  assign io_rf4debug_7 = rf_7; // @[RegisterFile.scala 46:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rf_1 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rf_2 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rf_3 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rf_4 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rf_5 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rf_6 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rf_7 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_write_0_rf_w) begin
      if (3'h1 == io_write_0_rd_addr) begin
        rf_1 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h2 == io_write_0_rd_addr) begin
        rf_2 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h3 == io_write_0_rd_addr) begin
        rf_3 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h4 == io_write_0_rd_addr) begin
        rf_4 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h5 == io_write_0_rd_addr) begin
        rf_5 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h6 == io_write_0_rd_addr) begin
        rf_6 <= io_write_0_data;
      end
    end
    if (io_write_0_rf_w) begin
      if (3'h7 == io_write_0_rd_addr) begin
        rf_7 <= io_write_0_data;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"we: %d, addr: %d, data: %d\n",io_write_0_rf_w,io_write_0_rd_addr,io_write_0_data); // @[RegisterFile.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"we: %d, addr: %d, data: %d\n",1'h0,3'h0,16'h0); // @[RegisterFile.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"rf: "); // @[RegisterFile.scala 52:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"0:%d, ",16'h0); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"1:%d, ",rf_1); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"2:%d, ",rf_2); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"3:%d, ",rf_3); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"4:%d, ",rf_4); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"5:%d, ",rf_5); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"6:%d, ",rf_6); // @[RegisterFile.scala 54:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"7:%d\n",rf_7); // @[RegisterFile.scala 55:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BusyBit(
  input        clock,
  input        reset,
  input        io_branch_mispredicted,
  input        io_branch_graduated,
  input  [2:0] io_release_0_rd_addr,
  input        io_release_0_rf_w,
  input  [2:0] io_req_rs_addr_0,
  input  [2:0] io_req_rs_addr_1,
  input        io_req_rd_w,
  input  [2:0] io_req_rd_addr,
  output       io_rs_available_0,
  output       io_rs_available_1
);
  reg  busy_bit_1; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_0;
  reg  busy_bit_2; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_1;
  reg  busy_bit_3; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_2;
  reg  busy_bit_4; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_3;
  reg  busy_bit_5; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_4;
  reg  busy_bit_6; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_5;
  reg  busy_bit_7; // @[BusyBit.scala 22:36]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[BusyBit.scala 26:78]
  wire  _T_2; // @[BusyBit.scala 26:65]
  wire  _GEN_784; // @[BusyBit.scala 27:27]
  wire  _GEN_1; // @[BusyBit.scala 27:27]
  wire  _GEN_2; // @[BusyBit.scala 27:27]
  wire  _GEN_3; // @[BusyBit.scala 27:27]
  wire  _GEN_4; // @[BusyBit.scala 27:27]
  wire  _GEN_5; // @[BusyBit.scala 27:27]
  wire  _GEN_6; // @[BusyBit.scala 27:27]
  wire  _GEN_7; // @[BusyBit.scala 27:27]
  wire  _T_7; // @[BusyBit.scala 27:27]
  wire  _T_9; // @[BusyBit.scala 26:78]
  wire  _T_10; // @[BusyBit.scala 26:65]
  wire  _GEN_785; // @[BusyBit.scala 27:27]
  wire  _GEN_9; // @[BusyBit.scala 27:27]
  wire  _GEN_10; // @[BusyBit.scala 27:27]
  wire  _GEN_11; // @[BusyBit.scala 27:27]
  wire  _GEN_12; // @[BusyBit.scala 27:27]
  wire  _GEN_13; // @[BusyBit.scala 27:27]
  wire  _GEN_14; // @[BusyBit.scala 27:27]
  wire  _GEN_15; // @[BusyBit.scala 27:27]
  wire  _T_15; // @[BusyBit.scala 27:27]
  wire  _T_17; // @[BusyBit.scala 31:30]
  wire  _GEN_17; // @[BusyBit.scala 32:39]
  wire  _GEN_18; // @[BusyBit.scala 32:39]
  wire  _GEN_19; // @[BusyBit.scala 32:39]
  wire  _GEN_20; // @[BusyBit.scala 32:39]
  wire  _GEN_21; // @[BusyBit.scala 32:39]
  wire  _GEN_22; // @[BusyBit.scala 32:39]
  wire  _GEN_23; // @[BusyBit.scala 32:39]
  wire  _T_18; // @[BusyBit.scala 33:62]
  wire  _T_19; // @[BusyBit.scala 33:37]
  wire  _T_20; // @[BusyBit.scala 35:48]
  wire  _T_21; // @[BusyBit.scala 35:30]
  wire  _GEN_786; // @[BusyBit.scala 36:32]
  wire  _GEN_33; // @[BusyBit.scala 36:32]
  wire  _GEN_787; // @[BusyBit.scala 36:32]
  wire  _GEN_34; // @[BusyBit.scala 36:32]
  wire  _GEN_788; // @[BusyBit.scala 36:32]
  wire  _GEN_35; // @[BusyBit.scala 36:32]
  wire  _GEN_789; // @[BusyBit.scala 36:32]
  wire  _GEN_36; // @[BusyBit.scala 36:32]
  wire  _GEN_790; // @[BusyBit.scala 36:32]
  wire  _GEN_37; // @[BusyBit.scala 36:32]
  wire  _GEN_791; // @[BusyBit.scala 36:32]
  wire  _GEN_38; // @[BusyBit.scala 36:32]
  wire  _GEN_792; // @[BusyBit.scala 36:32]
  wire  _GEN_39; // @[BusyBit.scala 36:32]
  wire  _GEN_41; // @[BusyBit.scala 35:57]
  wire  _GEN_42; // @[BusyBit.scala 35:57]
  wire  _GEN_43; // @[BusyBit.scala 35:57]
  wire  _GEN_44; // @[BusyBit.scala 35:57]
  wire  _GEN_45; // @[BusyBit.scala 35:57]
  wire  _GEN_46; // @[BusyBit.scala 35:57]
  wire  _GEN_47; // @[BusyBit.scala 35:57]
  wire  _GEN_49; // @[BusyBit.scala 33:71]
  wire  _GEN_50; // @[BusyBit.scala 33:71]
  wire  _GEN_51; // @[BusyBit.scala 33:71]
  wire  _GEN_52; // @[BusyBit.scala 33:71]
  wire  _GEN_53; // @[BusyBit.scala 33:71]
  wire  _GEN_54; // @[BusyBit.scala 33:71]
  wire  _GEN_55; // @[BusyBit.scala 33:71]
  wire  _GEN_57; // @[BusyBit.scala 31:57]
  wire  _GEN_58; // @[BusyBit.scala 31:57]
  wire  _GEN_59; // @[BusyBit.scala 31:57]
  wire  _GEN_60; // @[BusyBit.scala 31:57]
  wire  _GEN_61; // @[BusyBit.scala 31:57]
  wire  _GEN_62; // @[BusyBit.scala 31:57]
  wire  _GEN_63; // @[BusyBit.scala 31:57]
  wire  _GEN_65; // @[BusyBit.scala 32:39]
  wire  _GEN_66; // @[BusyBit.scala 32:39]
  wire  _GEN_67; // @[BusyBit.scala 32:39]
  wire  _GEN_68; // @[BusyBit.scala 32:39]
  wire  _GEN_69; // @[BusyBit.scala 32:39]
  wire  _GEN_70; // @[BusyBit.scala 32:39]
  wire  _GEN_71; // @[BusyBit.scala 32:39]
  wire  _T_23; // @[BusyBit.scala 33:62]
  wire  _T_24; // @[BusyBit.scala 33:37]
  wire  _T_25; // @[BusyBit.scala 35:48]
  wire  _T_26; // @[BusyBit.scala 35:30]
  wire  _GEN_81; // @[BusyBit.scala 36:32]
  wire  _GEN_82; // @[BusyBit.scala 36:32]
  wire  _GEN_83; // @[BusyBit.scala 36:32]
  wire  _GEN_84; // @[BusyBit.scala 36:32]
  wire  _GEN_85; // @[BusyBit.scala 36:32]
  wire  _GEN_86; // @[BusyBit.scala 36:32]
  wire  _GEN_87; // @[BusyBit.scala 36:32]
  wire  _GEN_89; // @[BusyBit.scala 35:57]
  wire  _GEN_90; // @[BusyBit.scala 35:57]
  wire  _GEN_91; // @[BusyBit.scala 35:57]
  wire  _GEN_92; // @[BusyBit.scala 35:57]
  wire  _GEN_93; // @[BusyBit.scala 35:57]
  wire  _GEN_94; // @[BusyBit.scala 35:57]
  wire  _GEN_95; // @[BusyBit.scala 35:57]
  wire  _GEN_97; // @[BusyBit.scala 33:71]
  wire  _GEN_98; // @[BusyBit.scala 33:71]
  wire  _GEN_99; // @[BusyBit.scala 33:71]
  wire  _GEN_100; // @[BusyBit.scala 33:71]
  wire  _GEN_101; // @[BusyBit.scala 33:71]
  wire  _GEN_102; // @[BusyBit.scala 33:71]
  wire  _GEN_103; // @[BusyBit.scala 33:71]
  wire  _GEN_105; // @[BusyBit.scala 31:57]
  wire  _GEN_106; // @[BusyBit.scala 31:57]
  wire  _GEN_107; // @[BusyBit.scala 31:57]
  wire  _GEN_108; // @[BusyBit.scala 31:57]
  wire  _GEN_109; // @[BusyBit.scala 31:57]
  wire  _GEN_110; // @[BusyBit.scala 31:57]
  wire  _GEN_111; // @[BusyBit.scala 31:57]
  wire  _GEN_113; // @[BusyBit.scala 32:39]
  wire  _GEN_114; // @[BusyBit.scala 32:39]
  wire  _GEN_115; // @[BusyBit.scala 32:39]
  wire  _GEN_116; // @[BusyBit.scala 32:39]
  wire  _GEN_117; // @[BusyBit.scala 32:39]
  wire  _GEN_118; // @[BusyBit.scala 32:39]
  wire  _GEN_119; // @[BusyBit.scala 32:39]
  wire  _T_28; // @[BusyBit.scala 33:62]
  wire  _T_29; // @[BusyBit.scala 33:37]
  wire  _T_30; // @[BusyBit.scala 35:48]
  wire  _T_31; // @[BusyBit.scala 35:30]
  wire  _GEN_129; // @[BusyBit.scala 36:32]
  wire  _GEN_130; // @[BusyBit.scala 36:32]
  wire  _GEN_131; // @[BusyBit.scala 36:32]
  wire  _GEN_132; // @[BusyBit.scala 36:32]
  wire  _GEN_133; // @[BusyBit.scala 36:32]
  wire  _GEN_134; // @[BusyBit.scala 36:32]
  wire  _GEN_135; // @[BusyBit.scala 36:32]
  wire  _GEN_137; // @[BusyBit.scala 35:57]
  wire  _GEN_138; // @[BusyBit.scala 35:57]
  wire  _GEN_139; // @[BusyBit.scala 35:57]
  wire  _GEN_140; // @[BusyBit.scala 35:57]
  wire  _GEN_141; // @[BusyBit.scala 35:57]
  wire  _GEN_142; // @[BusyBit.scala 35:57]
  wire  _GEN_143; // @[BusyBit.scala 35:57]
  wire  _GEN_145; // @[BusyBit.scala 33:71]
  wire  _GEN_146; // @[BusyBit.scala 33:71]
  wire  _GEN_147; // @[BusyBit.scala 33:71]
  wire  _GEN_148; // @[BusyBit.scala 33:71]
  wire  _GEN_149; // @[BusyBit.scala 33:71]
  wire  _GEN_150; // @[BusyBit.scala 33:71]
  wire  _GEN_151; // @[BusyBit.scala 33:71]
  wire  _GEN_153; // @[BusyBit.scala 31:57]
  wire  _GEN_154; // @[BusyBit.scala 31:57]
  wire  _GEN_155; // @[BusyBit.scala 31:57]
  wire  _GEN_156; // @[BusyBit.scala 31:57]
  wire  _GEN_157; // @[BusyBit.scala 31:57]
  wire  _GEN_158; // @[BusyBit.scala 31:57]
  wire  _GEN_159; // @[BusyBit.scala 31:57]
  wire  _GEN_161; // @[BusyBit.scala 32:39]
  wire  _GEN_162; // @[BusyBit.scala 32:39]
  wire  _GEN_163; // @[BusyBit.scala 32:39]
  wire  _GEN_164; // @[BusyBit.scala 32:39]
  wire  _GEN_165; // @[BusyBit.scala 32:39]
  wire  _GEN_166; // @[BusyBit.scala 32:39]
  wire  _GEN_167; // @[BusyBit.scala 32:39]
  wire  _T_33; // @[BusyBit.scala 33:62]
  wire  _T_34; // @[BusyBit.scala 33:37]
  wire  _T_35; // @[BusyBit.scala 35:48]
  wire  _T_36; // @[BusyBit.scala 35:30]
  wire  _GEN_177; // @[BusyBit.scala 36:32]
  wire  _GEN_178; // @[BusyBit.scala 36:32]
  wire  _GEN_179; // @[BusyBit.scala 36:32]
  wire  _GEN_180; // @[BusyBit.scala 36:32]
  wire  _GEN_181; // @[BusyBit.scala 36:32]
  wire  _GEN_182; // @[BusyBit.scala 36:32]
  wire  _GEN_183; // @[BusyBit.scala 36:32]
  wire  _GEN_185; // @[BusyBit.scala 35:57]
  wire  _GEN_186; // @[BusyBit.scala 35:57]
  wire  _GEN_187; // @[BusyBit.scala 35:57]
  wire  _GEN_188; // @[BusyBit.scala 35:57]
  wire  _GEN_189; // @[BusyBit.scala 35:57]
  wire  _GEN_190; // @[BusyBit.scala 35:57]
  wire  _GEN_191; // @[BusyBit.scala 35:57]
  wire  _GEN_193; // @[BusyBit.scala 33:71]
  wire  _GEN_194; // @[BusyBit.scala 33:71]
  wire  _GEN_195; // @[BusyBit.scala 33:71]
  wire  _GEN_196; // @[BusyBit.scala 33:71]
  wire  _GEN_197; // @[BusyBit.scala 33:71]
  wire  _GEN_198; // @[BusyBit.scala 33:71]
  wire  _GEN_199; // @[BusyBit.scala 33:71]
  wire  _GEN_201; // @[BusyBit.scala 31:57]
  wire  _GEN_202; // @[BusyBit.scala 31:57]
  wire  _GEN_203; // @[BusyBit.scala 31:57]
  wire  _GEN_204; // @[BusyBit.scala 31:57]
  wire  _GEN_205; // @[BusyBit.scala 31:57]
  wire  _GEN_206; // @[BusyBit.scala 31:57]
  wire  _GEN_207; // @[BusyBit.scala 31:57]
  wire  _GEN_209; // @[BusyBit.scala 32:39]
  wire  _GEN_210; // @[BusyBit.scala 32:39]
  wire  _GEN_211; // @[BusyBit.scala 32:39]
  wire  _GEN_212; // @[BusyBit.scala 32:39]
  wire  _GEN_213; // @[BusyBit.scala 32:39]
  wire  _GEN_214; // @[BusyBit.scala 32:39]
  wire  _GEN_215; // @[BusyBit.scala 32:39]
  wire  _T_38; // @[BusyBit.scala 33:62]
  wire  _T_39; // @[BusyBit.scala 33:37]
  wire  _T_40; // @[BusyBit.scala 35:48]
  wire  _T_41; // @[BusyBit.scala 35:30]
  wire  _GEN_225; // @[BusyBit.scala 36:32]
  wire  _GEN_226; // @[BusyBit.scala 36:32]
  wire  _GEN_227; // @[BusyBit.scala 36:32]
  wire  _GEN_228; // @[BusyBit.scala 36:32]
  wire  _GEN_229; // @[BusyBit.scala 36:32]
  wire  _GEN_230; // @[BusyBit.scala 36:32]
  wire  _GEN_231; // @[BusyBit.scala 36:32]
  wire  _GEN_233; // @[BusyBit.scala 35:57]
  wire  _GEN_234; // @[BusyBit.scala 35:57]
  wire  _GEN_235; // @[BusyBit.scala 35:57]
  wire  _GEN_236; // @[BusyBit.scala 35:57]
  wire  _GEN_237; // @[BusyBit.scala 35:57]
  wire  _GEN_238; // @[BusyBit.scala 35:57]
  wire  _GEN_239; // @[BusyBit.scala 35:57]
  wire  _GEN_241; // @[BusyBit.scala 33:71]
  wire  _GEN_242; // @[BusyBit.scala 33:71]
  wire  _GEN_243; // @[BusyBit.scala 33:71]
  wire  _GEN_244; // @[BusyBit.scala 33:71]
  wire  _GEN_245; // @[BusyBit.scala 33:71]
  wire  _GEN_246; // @[BusyBit.scala 33:71]
  wire  _GEN_247; // @[BusyBit.scala 33:71]
  wire  _GEN_249; // @[BusyBit.scala 31:57]
  wire  _GEN_250; // @[BusyBit.scala 31:57]
  wire  _GEN_251; // @[BusyBit.scala 31:57]
  wire  _GEN_252; // @[BusyBit.scala 31:57]
  wire  _GEN_253; // @[BusyBit.scala 31:57]
  wire  _GEN_254; // @[BusyBit.scala 31:57]
  wire  _GEN_255; // @[BusyBit.scala 31:57]
  wire  _GEN_257; // @[BusyBit.scala 32:39]
  wire  _GEN_258; // @[BusyBit.scala 32:39]
  wire  _GEN_259; // @[BusyBit.scala 32:39]
  wire  _GEN_260; // @[BusyBit.scala 32:39]
  wire  _GEN_261; // @[BusyBit.scala 32:39]
  wire  _GEN_262; // @[BusyBit.scala 32:39]
  wire  _GEN_263; // @[BusyBit.scala 32:39]
  wire  _T_43; // @[BusyBit.scala 33:62]
  wire  _T_44; // @[BusyBit.scala 33:37]
  wire  _T_45; // @[BusyBit.scala 35:48]
  wire  _T_46; // @[BusyBit.scala 35:30]
  wire  _GEN_273; // @[BusyBit.scala 36:32]
  wire  _GEN_274; // @[BusyBit.scala 36:32]
  wire  _GEN_275; // @[BusyBit.scala 36:32]
  wire  _GEN_276; // @[BusyBit.scala 36:32]
  wire  _GEN_277; // @[BusyBit.scala 36:32]
  wire  _GEN_278; // @[BusyBit.scala 36:32]
  wire  _GEN_279; // @[BusyBit.scala 36:32]
  wire  _GEN_281; // @[BusyBit.scala 35:57]
  wire  _GEN_282; // @[BusyBit.scala 35:57]
  wire  _GEN_283; // @[BusyBit.scala 35:57]
  wire  _GEN_284; // @[BusyBit.scala 35:57]
  wire  _GEN_285; // @[BusyBit.scala 35:57]
  wire  _GEN_286; // @[BusyBit.scala 35:57]
  wire  _GEN_287; // @[BusyBit.scala 35:57]
  wire  _GEN_289; // @[BusyBit.scala 33:71]
  wire  _GEN_290; // @[BusyBit.scala 33:71]
  wire  _GEN_291; // @[BusyBit.scala 33:71]
  wire  _GEN_292; // @[BusyBit.scala 33:71]
  wire  _GEN_293; // @[BusyBit.scala 33:71]
  wire  _GEN_294; // @[BusyBit.scala 33:71]
  wire  _GEN_295; // @[BusyBit.scala 33:71]
  wire  _GEN_297; // @[BusyBit.scala 31:57]
  wire  _GEN_298; // @[BusyBit.scala 31:57]
  wire  _GEN_299; // @[BusyBit.scala 31:57]
  wire  _GEN_300; // @[BusyBit.scala 31:57]
  wire  _GEN_301; // @[BusyBit.scala 31:57]
  wire  _GEN_302; // @[BusyBit.scala 31:57]
  wire  _GEN_303; // @[BusyBit.scala 31:57]
  wire  _GEN_305; // @[BusyBit.scala 32:39]
  wire  _GEN_306; // @[BusyBit.scala 32:39]
  wire  _GEN_307; // @[BusyBit.scala 32:39]
  wire  _GEN_308; // @[BusyBit.scala 32:39]
  wire  _GEN_309; // @[BusyBit.scala 32:39]
  wire  _GEN_310; // @[BusyBit.scala 32:39]
  wire  _GEN_311; // @[BusyBit.scala 32:39]
  wire  _T_48; // @[BusyBit.scala 33:62]
  wire  _T_49; // @[BusyBit.scala 33:37]
  wire  _T_50; // @[BusyBit.scala 35:48]
  wire  _T_51; // @[BusyBit.scala 35:30]
  wire  _GEN_321; // @[BusyBit.scala 36:32]
  wire  _GEN_322; // @[BusyBit.scala 36:32]
  wire  _GEN_323; // @[BusyBit.scala 36:32]
  wire  _GEN_324; // @[BusyBit.scala 36:32]
  wire  _GEN_325; // @[BusyBit.scala 36:32]
  wire  _GEN_326; // @[BusyBit.scala 36:32]
  wire  _GEN_327; // @[BusyBit.scala 36:32]
  wire  _GEN_329; // @[BusyBit.scala 35:57]
  wire  _GEN_330; // @[BusyBit.scala 35:57]
  wire  _GEN_331; // @[BusyBit.scala 35:57]
  wire  _GEN_332; // @[BusyBit.scala 35:57]
  wire  _GEN_333; // @[BusyBit.scala 35:57]
  wire  _GEN_334; // @[BusyBit.scala 35:57]
  wire  _GEN_335; // @[BusyBit.scala 35:57]
  wire  _GEN_337; // @[BusyBit.scala 33:71]
  wire  _GEN_338; // @[BusyBit.scala 33:71]
  wire  _GEN_339; // @[BusyBit.scala 33:71]
  wire  _GEN_340; // @[BusyBit.scala 33:71]
  wire  _GEN_341; // @[BusyBit.scala 33:71]
  wire  _GEN_342; // @[BusyBit.scala 33:71]
  wire  _GEN_343; // @[BusyBit.scala 33:71]
  wire  _GEN_345; // @[BusyBit.scala 31:57]
  wire  _GEN_346; // @[BusyBit.scala 31:57]
  wire  _GEN_347; // @[BusyBit.scala 31:57]
  wire  _GEN_348; // @[BusyBit.scala 31:57]
  wire  _GEN_349; // @[BusyBit.scala 31:57]
  wire  _GEN_350; // @[BusyBit.scala 31:57]
  wire  _GEN_351; // @[BusyBit.scala 31:57]
  wire  _GEN_353; // @[BusyBit.scala 32:39]
  wire  _GEN_354; // @[BusyBit.scala 32:39]
  wire  _GEN_355; // @[BusyBit.scala 32:39]
  wire  _GEN_356; // @[BusyBit.scala 32:39]
  wire  _GEN_357; // @[BusyBit.scala 32:39]
  wire  _GEN_358; // @[BusyBit.scala 32:39]
  wire  _GEN_359; // @[BusyBit.scala 32:39]
  wire  _T_53; // @[BusyBit.scala 33:62]
  wire  _T_54; // @[BusyBit.scala 33:37]
  wire  _T_55; // @[BusyBit.scala 35:48]
  wire  _T_56; // @[BusyBit.scala 35:30]
  wire  _GEN_369; // @[BusyBit.scala 36:32]
  wire  _GEN_370; // @[BusyBit.scala 36:32]
  wire  _GEN_371; // @[BusyBit.scala 36:32]
  wire  _GEN_372; // @[BusyBit.scala 36:32]
  wire  _GEN_373; // @[BusyBit.scala 36:32]
  wire  _GEN_374; // @[BusyBit.scala 36:32]
  wire  _GEN_375; // @[BusyBit.scala 36:32]
  wire  _GEN_377; // @[BusyBit.scala 35:57]
  wire  _GEN_378; // @[BusyBit.scala 35:57]
  wire  _GEN_379; // @[BusyBit.scala 35:57]
  wire  _GEN_380; // @[BusyBit.scala 35:57]
  wire  _GEN_381; // @[BusyBit.scala 35:57]
  wire  _GEN_382; // @[BusyBit.scala 35:57]
  wire  _GEN_383; // @[BusyBit.scala 35:57]
  wire  _GEN_385; // @[BusyBit.scala 33:71]
  wire  _GEN_386; // @[BusyBit.scala 33:71]
  wire  _GEN_387; // @[BusyBit.scala 33:71]
  wire  _GEN_388; // @[BusyBit.scala 33:71]
  wire  _GEN_389; // @[BusyBit.scala 33:71]
  wire  _GEN_390; // @[BusyBit.scala 33:71]
  wire  _GEN_391; // @[BusyBit.scala 33:71]
  wire  _GEN_393; // @[BusyBit.scala 31:57]
  wire  _GEN_394; // @[BusyBit.scala 31:57]
  wire  _GEN_395; // @[BusyBit.scala 31:57]
  wire  _GEN_396; // @[BusyBit.scala 31:57]
  wire  _GEN_397; // @[BusyBit.scala 31:57]
  wire  _GEN_398; // @[BusyBit.scala 31:57]
  wire  _GEN_399; // @[BusyBit.scala 31:57]
  wire  _GEN_417; // @[BusyBit.scala 36:32]
  wire  _GEN_418; // @[BusyBit.scala 36:32]
  wire  _GEN_419; // @[BusyBit.scala 36:32]
  wire  _GEN_420; // @[BusyBit.scala 36:32]
  wire  _GEN_421; // @[BusyBit.scala 36:32]
  wire  _GEN_422; // @[BusyBit.scala 36:32]
  wire  _GEN_423; // @[BusyBit.scala 36:32]
  wire  _GEN_425; // @[BusyBit.scala 35:57]
  wire  _GEN_426; // @[BusyBit.scala 35:57]
  wire  _GEN_427; // @[BusyBit.scala 35:57]
  wire  _GEN_428; // @[BusyBit.scala 35:57]
  wire  _GEN_429; // @[BusyBit.scala 35:57]
  wire  _GEN_430; // @[BusyBit.scala 35:57]
  wire  _GEN_431; // @[BusyBit.scala 35:57]
  wire  _GEN_441; // @[BusyBit.scala 31:57]
  wire  _GEN_442; // @[BusyBit.scala 31:57]
  wire  _GEN_443; // @[BusyBit.scala 31:57]
  wire  _GEN_444; // @[BusyBit.scala 31:57]
  wire  _GEN_445; // @[BusyBit.scala 31:57]
  wire  _GEN_446; // @[BusyBit.scala 31:57]
  wire  _GEN_447; // @[BusyBit.scala 31:57]
  wire  _GEN_465; // @[BusyBit.scala 36:32]
  wire  _GEN_466; // @[BusyBit.scala 36:32]
  wire  _GEN_467; // @[BusyBit.scala 36:32]
  wire  _GEN_468; // @[BusyBit.scala 36:32]
  wire  _GEN_469; // @[BusyBit.scala 36:32]
  wire  _GEN_470; // @[BusyBit.scala 36:32]
  wire  _GEN_471; // @[BusyBit.scala 36:32]
  wire  _GEN_473; // @[BusyBit.scala 35:57]
  wire  _GEN_474; // @[BusyBit.scala 35:57]
  wire  _GEN_475; // @[BusyBit.scala 35:57]
  wire  _GEN_476; // @[BusyBit.scala 35:57]
  wire  _GEN_477; // @[BusyBit.scala 35:57]
  wire  _GEN_478; // @[BusyBit.scala 35:57]
  wire  _GEN_479; // @[BusyBit.scala 35:57]
  wire  _GEN_489; // @[BusyBit.scala 31:57]
  wire  _GEN_490; // @[BusyBit.scala 31:57]
  wire  _GEN_491; // @[BusyBit.scala 31:57]
  wire  _GEN_492; // @[BusyBit.scala 31:57]
  wire  _GEN_493; // @[BusyBit.scala 31:57]
  wire  _GEN_494; // @[BusyBit.scala 31:57]
  wire  _GEN_495; // @[BusyBit.scala 31:57]
  wire  _GEN_513; // @[BusyBit.scala 36:32]
  wire  _GEN_514; // @[BusyBit.scala 36:32]
  wire  _GEN_515; // @[BusyBit.scala 36:32]
  wire  _GEN_516; // @[BusyBit.scala 36:32]
  wire  _GEN_517; // @[BusyBit.scala 36:32]
  wire  _GEN_518; // @[BusyBit.scala 36:32]
  wire  _GEN_519; // @[BusyBit.scala 36:32]
  wire  _GEN_521; // @[BusyBit.scala 35:57]
  wire  _GEN_522; // @[BusyBit.scala 35:57]
  wire  _GEN_523; // @[BusyBit.scala 35:57]
  wire  _GEN_524; // @[BusyBit.scala 35:57]
  wire  _GEN_525; // @[BusyBit.scala 35:57]
  wire  _GEN_526; // @[BusyBit.scala 35:57]
  wire  _GEN_527; // @[BusyBit.scala 35:57]
  wire  _GEN_537; // @[BusyBit.scala 31:57]
  wire  _GEN_538; // @[BusyBit.scala 31:57]
  wire  _GEN_539; // @[BusyBit.scala 31:57]
  wire  _GEN_540; // @[BusyBit.scala 31:57]
  wire  _GEN_541; // @[BusyBit.scala 31:57]
  wire  _GEN_542; // @[BusyBit.scala 31:57]
  wire  _GEN_543; // @[BusyBit.scala 31:57]
  wire  _GEN_561; // @[BusyBit.scala 36:32]
  wire  _GEN_562; // @[BusyBit.scala 36:32]
  wire  _GEN_563; // @[BusyBit.scala 36:32]
  wire  _GEN_564; // @[BusyBit.scala 36:32]
  wire  _GEN_565; // @[BusyBit.scala 36:32]
  wire  _GEN_566; // @[BusyBit.scala 36:32]
  wire  _GEN_567; // @[BusyBit.scala 36:32]
  wire  _GEN_569; // @[BusyBit.scala 35:57]
  wire  _GEN_570; // @[BusyBit.scala 35:57]
  wire  _GEN_571; // @[BusyBit.scala 35:57]
  wire  _GEN_572; // @[BusyBit.scala 35:57]
  wire  _GEN_573; // @[BusyBit.scala 35:57]
  wire  _GEN_574; // @[BusyBit.scala 35:57]
  wire  _GEN_575; // @[BusyBit.scala 35:57]
  wire  _GEN_585; // @[BusyBit.scala 31:57]
  wire  _GEN_586; // @[BusyBit.scala 31:57]
  wire  _GEN_587; // @[BusyBit.scala 31:57]
  wire  _GEN_588; // @[BusyBit.scala 31:57]
  wire  _GEN_589; // @[BusyBit.scala 31:57]
  wire  _GEN_590; // @[BusyBit.scala 31:57]
  wire  _GEN_591; // @[BusyBit.scala 31:57]
  wire  _GEN_609; // @[BusyBit.scala 36:32]
  wire  _GEN_610; // @[BusyBit.scala 36:32]
  wire  _GEN_611; // @[BusyBit.scala 36:32]
  wire  _GEN_612; // @[BusyBit.scala 36:32]
  wire  _GEN_613; // @[BusyBit.scala 36:32]
  wire  _GEN_614; // @[BusyBit.scala 36:32]
  wire  _GEN_615; // @[BusyBit.scala 36:32]
  wire  _GEN_617; // @[BusyBit.scala 35:57]
  wire  _GEN_618; // @[BusyBit.scala 35:57]
  wire  _GEN_619; // @[BusyBit.scala 35:57]
  wire  _GEN_620; // @[BusyBit.scala 35:57]
  wire  _GEN_621; // @[BusyBit.scala 35:57]
  wire  _GEN_622; // @[BusyBit.scala 35:57]
  wire  _GEN_623; // @[BusyBit.scala 35:57]
  wire  _GEN_633; // @[BusyBit.scala 31:57]
  wire  _GEN_634; // @[BusyBit.scala 31:57]
  wire  _GEN_635; // @[BusyBit.scala 31:57]
  wire  _GEN_636; // @[BusyBit.scala 31:57]
  wire  _GEN_637; // @[BusyBit.scala 31:57]
  wire  _GEN_638; // @[BusyBit.scala 31:57]
  wire  _GEN_639; // @[BusyBit.scala 31:57]
  wire  _GEN_657; // @[BusyBit.scala 36:32]
  wire  _GEN_658; // @[BusyBit.scala 36:32]
  wire  _GEN_659; // @[BusyBit.scala 36:32]
  wire  _GEN_660; // @[BusyBit.scala 36:32]
  wire  _GEN_661; // @[BusyBit.scala 36:32]
  wire  _GEN_662; // @[BusyBit.scala 36:32]
  wire  _GEN_663; // @[BusyBit.scala 36:32]
  wire  _GEN_665; // @[BusyBit.scala 35:57]
  wire  _GEN_666; // @[BusyBit.scala 35:57]
  wire  _GEN_667; // @[BusyBit.scala 35:57]
  wire  _GEN_668; // @[BusyBit.scala 35:57]
  wire  _GEN_669; // @[BusyBit.scala 35:57]
  wire  _GEN_670; // @[BusyBit.scala 35:57]
  wire  _GEN_671; // @[BusyBit.scala 35:57]
  wire  _GEN_681; // @[BusyBit.scala 31:57]
  wire  _GEN_682; // @[BusyBit.scala 31:57]
  wire  _GEN_683; // @[BusyBit.scala 31:57]
  wire  _GEN_684; // @[BusyBit.scala 31:57]
  wire  _GEN_685; // @[BusyBit.scala 31:57]
  wire  _GEN_686; // @[BusyBit.scala 31:57]
  wire  _GEN_687; // @[BusyBit.scala 31:57]
  wire  _GEN_705; // @[BusyBit.scala 36:32]
  wire  _GEN_706; // @[BusyBit.scala 36:32]
  wire  _GEN_707; // @[BusyBit.scala 36:32]
  wire  _GEN_708; // @[BusyBit.scala 36:32]
  wire  _GEN_709; // @[BusyBit.scala 36:32]
  wire  _GEN_710; // @[BusyBit.scala 36:32]
  wire  _GEN_711; // @[BusyBit.scala 36:32]
  wire  _GEN_713; // @[BusyBit.scala 35:57]
  wire  _GEN_714; // @[BusyBit.scala 35:57]
  wire  _GEN_715; // @[BusyBit.scala 35:57]
  wire  _GEN_716; // @[BusyBit.scala 35:57]
  wire  _GEN_717; // @[BusyBit.scala 35:57]
  wire  _GEN_718; // @[BusyBit.scala 35:57]
  wire  _GEN_719; // @[BusyBit.scala 35:57]
  wire  _GEN_729; // @[BusyBit.scala 31:57]
  wire  _GEN_730; // @[BusyBit.scala 31:57]
  wire  _GEN_731; // @[BusyBit.scala 31:57]
  wire  _GEN_732; // @[BusyBit.scala 31:57]
  wire  _GEN_733; // @[BusyBit.scala 31:57]
  wire  _GEN_734; // @[BusyBit.scala 31:57]
  wire  _GEN_735; // @[BusyBit.scala 31:57]
  wire  _GEN_753; // @[BusyBit.scala 36:32]
  wire  _GEN_754; // @[BusyBit.scala 36:32]
  wire  _GEN_755; // @[BusyBit.scala 36:32]
  wire  _GEN_756; // @[BusyBit.scala 36:32]
  wire  _GEN_757; // @[BusyBit.scala 36:32]
  wire  _GEN_758; // @[BusyBit.scala 36:32]
  wire  _GEN_759; // @[BusyBit.scala 36:32]
  wire  _T_97; // @[BusyBit.scala 40:9]
  wire  _T_98; // @[BusyBit.scala 40:9]
  assign _T_1 = io_release_0_rd_addr == io_req_rs_addr_0; // @[BusyBit.scala 26:78]
  assign _T_2 = io_release_0_rf_w & _T_1; // @[BusyBit.scala 26:65]
  assign _GEN_784 = 3'h1 == io_req_rs_addr_0; // @[BusyBit.scala 27:27]
  assign _GEN_1 = _GEN_784 & busy_bit_1; // @[BusyBit.scala 27:27]
  assign _GEN_2 = 3'h2 == io_req_rs_addr_0 ? busy_bit_2 : _GEN_1; // @[BusyBit.scala 27:27]
  assign _GEN_3 = 3'h3 == io_req_rs_addr_0 ? busy_bit_3 : _GEN_2; // @[BusyBit.scala 27:27]
  assign _GEN_4 = 3'h4 == io_req_rs_addr_0 ? busy_bit_4 : _GEN_3; // @[BusyBit.scala 27:27]
  assign _GEN_5 = 3'h5 == io_req_rs_addr_0 ? busy_bit_5 : _GEN_4; // @[BusyBit.scala 27:27]
  assign _GEN_6 = 3'h6 == io_req_rs_addr_0 ? busy_bit_6 : _GEN_5; // @[BusyBit.scala 27:27]
  assign _GEN_7 = 3'h7 == io_req_rs_addr_0 ? busy_bit_7 : _GEN_6; // @[BusyBit.scala 27:27]
  assign _T_7 = _GEN_7 == 1'h0; // @[BusyBit.scala 27:27]
  assign _T_9 = io_release_0_rd_addr == io_req_rs_addr_1; // @[BusyBit.scala 26:78]
  assign _T_10 = io_release_0_rf_w & _T_9; // @[BusyBit.scala 26:65]
  assign _GEN_785 = 3'h1 == io_req_rs_addr_1; // @[BusyBit.scala 27:27]
  assign _GEN_9 = _GEN_785 & busy_bit_1; // @[BusyBit.scala 27:27]
  assign _GEN_10 = 3'h2 == io_req_rs_addr_1 ? busy_bit_2 : _GEN_9; // @[BusyBit.scala 27:27]
  assign _GEN_11 = 3'h3 == io_req_rs_addr_1 ? busy_bit_3 : _GEN_10; // @[BusyBit.scala 27:27]
  assign _GEN_12 = 3'h4 == io_req_rs_addr_1 ? busy_bit_4 : _GEN_11; // @[BusyBit.scala 27:27]
  assign _GEN_13 = 3'h5 == io_req_rs_addr_1 ? busy_bit_5 : _GEN_12; // @[BusyBit.scala 27:27]
  assign _GEN_14 = 3'h6 == io_req_rs_addr_1 ? busy_bit_6 : _GEN_13; // @[BusyBit.scala 27:27]
  assign _GEN_15 = 3'h7 == io_req_rs_addr_1 ? busy_bit_7 : _GEN_14; // @[BusyBit.scala 27:27]
  assign _T_15 = _GEN_15 == 1'h0; // @[BusyBit.scala 27:27]
  assign _T_17 = io_branch_graduated & io_branch_mispredicted; // @[BusyBit.scala 31:30]
  assign _GEN_17 = 3'h1 == io_release_0_rd_addr ? 1'h0 : busy_bit_1; // @[BusyBit.scala 32:39]
  assign _GEN_18 = 3'h2 == io_release_0_rd_addr ? 1'h0 : busy_bit_2; // @[BusyBit.scala 32:39]
  assign _GEN_19 = 3'h3 == io_release_0_rd_addr ? 1'h0 : busy_bit_3; // @[BusyBit.scala 32:39]
  assign _GEN_20 = 3'h4 == io_release_0_rd_addr ? 1'h0 : busy_bit_4; // @[BusyBit.scala 32:39]
  assign _GEN_21 = 3'h5 == io_release_0_rd_addr ? 1'h0 : busy_bit_5; // @[BusyBit.scala 32:39]
  assign _GEN_22 = 3'h6 == io_release_0_rd_addr ? 1'h0 : busy_bit_6; // @[BusyBit.scala 32:39]
  assign _GEN_23 = 3'h7 == io_release_0_rd_addr ? 1'h0 : busy_bit_7; // @[BusyBit.scala 32:39]
  assign _T_18 = io_release_0_rd_addr == 3'h0; // @[BusyBit.scala 33:62]
  assign _T_19 = io_release_0_rf_w & _T_18; // @[BusyBit.scala 33:37]
  assign _T_20 = io_req_rd_addr == 3'h0; // @[BusyBit.scala 35:48]
  assign _T_21 = io_req_rd_w & _T_20; // @[BusyBit.scala 35:30]
  assign _GEN_786 = 3'h1 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_33 = _GEN_786 | busy_bit_1; // @[BusyBit.scala 36:32]
  assign _GEN_787 = 3'h2 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_34 = _GEN_787 | busy_bit_2; // @[BusyBit.scala 36:32]
  assign _GEN_788 = 3'h3 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_35 = _GEN_788 | busy_bit_3; // @[BusyBit.scala 36:32]
  assign _GEN_789 = 3'h4 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_36 = _GEN_789 | busy_bit_4; // @[BusyBit.scala 36:32]
  assign _GEN_790 = 3'h5 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_37 = _GEN_790 | busy_bit_5; // @[BusyBit.scala 36:32]
  assign _GEN_791 = 3'h6 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_38 = _GEN_791 | busy_bit_6; // @[BusyBit.scala 36:32]
  assign _GEN_792 = 3'h7 == io_req_rd_addr; // @[BusyBit.scala 36:32]
  assign _GEN_39 = _GEN_792 | busy_bit_7; // @[BusyBit.scala 36:32]
  assign _GEN_41 = _T_21 ? _GEN_33 : busy_bit_1; // @[BusyBit.scala 35:57]
  assign _GEN_42 = _T_21 ? _GEN_34 : busy_bit_2; // @[BusyBit.scala 35:57]
  assign _GEN_43 = _T_21 ? _GEN_35 : busy_bit_3; // @[BusyBit.scala 35:57]
  assign _GEN_44 = _T_21 ? _GEN_36 : busy_bit_4; // @[BusyBit.scala 35:57]
  assign _GEN_45 = _T_21 ? _GEN_37 : busy_bit_5; // @[BusyBit.scala 35:57]
  assign _GEN_46 = _T_21 ? _GEN_38 : busy_bit_6; // @[BusyBit.scala 35:57]
  assign _GEN_47 = _T_21 ? _GEN_39 : busy_bit_7; // @[BusyBit.scala 35:57]
  assign _GEN_49 = _T_19 ? _GEN_17 : _GEN_41; // @[BusyBit.scala 33:71]
  assign _GEN_50 = _T_19 ? _GEN_18 : _GEN_42; // @[BusyBit.scala 33:71]
  assign _GEN_51 = _T_19 ? _GEN_19 : _GEN_43; // @[BusyBit.scala 33:71]
  assign _GEN_52 = _T_19 ? _GEN_20 : _GEN_44; // @[BusyBit.scala 33:71]
  assign _GEN_53 = _T_19 ? _GEN_21 : _GEN_45; // @[BusyBit.scala 33:71]
  assign _GEN_54 = _T_19 ? _GEN_22 : _GEN_46; // @[BusyBit.scala 33:71]
  assign _GEN_55 = _T_19 ? _GEN_23 : _GEN_47; // @[BusyBit.scala 33:71]
  assign _GEN_57 = _T_17 ? _GEN_17 : _GEN_49; // @[BusyBit.scala 31:57]
  assign _GEN_58 = _T_17 ? _GEN_18 : _GEN_50; // @[BusyBit.scala 31:57]
  assign _GEN_59 = _T_17 ? _GEN_19 : _GEN_51; // @[BusyBit.scala 31:57]
  assign _GEN_60 = _T_17 ? _GEN_20 : _GEN_52; // @[BusyBit.scala 31:57]
  assign _GEN_61 = _T_17 ? _GEN_21 : _GEN_53; // @[BusyBit.scala 31:57]
  assign _GEN_62 = _T_17 ? _GEN_22 : _GEN_54; // @[BusyBit.scala 31:57]
  assign _GEN_63 = _T_17 ? _GEN_23 : _GEN_55; // @[BusyBit.scala 31:57]
  assign _GEN_65 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_57; // @[BusyBit.scala 32:39]
  assign _GEN_66 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_58; // @[BusyBit.scala 32:39]
  assign _GEN_67 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_59; // @[BusyBit.scala 32:39]
  assign _GEN_68 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_60; // @[BusyBit.scala 32:39]
  assign _GEN_69 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_61; // @[BusyBit.scala 32:39]
  assign _GEN_70 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_62; // @[BusyBit.scala 32:39]
  assign _GEN_71 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_63; // @[BusyBit.scala 32:39]
  assign _T_23 = io_release_0_rd_addr == 3'h1; // @[BusyBit.scala 33:62]
  assign _T_24 = io_release_0_rf_w & _T_23; // @[BusyBit.scala 33:37]
  assign _T_25 = io_req_rd_addr == 3'h1; // @[BusyBit.scala 35:48]
  assign _T_26 = io_req_rd_w & _T_25; // @[BusyBit.scala 35:30]
  assign _GEN_81 = _GEN_786 | _GEN_57; // @[BusyBit.scala 36:32]
  assign _GEN_82 = _GEN_787 | _GEN_58; // @[BusyBit.scala 36:32]
  assign _GEN_83 = _GEN_788 | _GEN_59; // @[BusyBit.scala 36:32]
  assign _GEN_84 = _GEN_789 | _GEN_60; // @[BusyBit.scala 36:32]
  assign _GEN_85 = _GEN_790 | _GEN_61; // @[BusyBit.scala 36:32]
  assign _GEN_86 = _GEN_791 | _GEN_62; // @[BusyBit.scala 36:32]
  assign _GEN_87 = _GEN_792 | _GEN_63; // @[BusyBit.scala 36:32]
  assign _GEN_89 = _T_26 ? _GEN_81 : _GEN_57; // @[BusyBit.scala 35:57]
  assign _GEN_90 = _T_26 ? _GEN_82 : _GEN_58; // @[BusyBit.scala 35:57]
  assign _GEN_91 = _T_26 ? _GEN_83 : _GEN_59; // @[BusyBit.scala 35:57]
  assign _GEN_92 = _T_26 ? _GEN_84 : _GEN_60; // @[BusyBit.scala 35:57]
  assign _GEN_93 = _T_26 ? _GEN_85 : _GEN_61; // @[BusyBit.scala 35:57]
  assign _GEN_94 = _T_26 ? _GEN_86 : _GEN_62; // @[BusyBit.scala 35:57]
  assign _GEN_95 = _T_26 ? _GEN_87 : _GEN_63; // @[BusyBit.scala 35:57]
  assign _GEN_97 = _T_24 ? _GEN_65 : _GEN_89; // @[BusyBit.scala 33:71]
  assign _GEN_98 = _T_24 ? _GEN_66 : _GEN_90; // @[BusyBit.scala 33:71]
  assign _GEN_99 = _T_24 ? _GEN_67 : _GEN_91; // @[BusyBit.scala 33:71]
  assign _GEN_100 = _T_24 ? _GEN_68 : _GEN_92; // @[BusyBit.scala 33:71]
  assign _GEN_101 = _T_24 ? _GEN_69 : _GEN_93; // @[BusyBit.scala 33:71]
  assign _GEN_102 = _T_24 ? _GEN_70 : _GEN_94; // @[BusyBit.scala 33:71]
  assign _GEN_103 = _T_24 ? _GEN_71 : _GEN_95; // @[BusyBit.scala 33:71]
  assign _GEN_105 = _T_17 ? _GEN_65 : _GEN_97; // @[BusyBit.scala 31:57]
  assign _GEN_106 = _T_17 ? _GEN_66 : _GEN_98; // @[BusyBit.scala 31:57]
  assign _GEN_107 = _T_17 ? _GEN_67 : _GEN_99; // @[BusyBit.scala 31:57]
  assign _GEN_108 = _T_17 ? _GEN_68 : _GEN_100; // @[BusyBit.scala 31:57]
  assign _GEN_109 = _T_17 ? _GEN_69 : _GEN_101; // @[BusyBit.scala 31:57]
  assign _GEN_110 = _T_17 ? _GEN_70 : _GEN_102; // @[BusyBit.scala 31:57]
  assign _GEN_111 = _T_17 ? _GEN_71 : _GEN_103; // @[BusyBit.scala 31:57]
  assign _GEN_113 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_105; // @[BusyBit.scala 32:39]
  assign _GEN_114 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_106; // @[BusyBit.scala 32:39]
  assign _GEN_115 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_107; // @[BusyBit.scala 32:39]
  assign _GEN_116 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_108; // @[BusyBit.scala 32:39]
  assign _GEN_117 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_109; // @[BusyBit.scala 32:39]
  assign _GEN_118 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_110; // @[BusyBit.scala 32:39]
  assign _GEN_119 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_111; // @[BusyBit.scala 32:39]
  assign _T_28 = io_release_0_rd_addr == 3'h2; // @[BusyBit.scala 33:62]
  assign _T_29 = io_release_0_rf_w & _T_28; // @[BusyBit.scala 33:37]
  assign _T_30 = io_req_rd_addr == 3'h2; // @[BusyBit.scala 35:48]
  assign _T_31 = io_req_rd_w & _T_30; // @[BusyBit.scala 35:30]
  assign _GEN_129 = _GEN_786 | _GEN_105; // @[BusyBit.scala 36:32]
  assign _GEN_130 = _GEN_787 | _GEN_106; // @[BusyBit.scala 36:32]
  assign _GEN_131 = _GEN_788 | _GEN_107; // @[BusyBit.scala 36:32]
  assign _GEN_132 = _GEN_789 | _GEN_108; // @[BusyBit.scala 36:32]
  assign _GEN_133 = _GEN_790 | _GEN_109; // @[BusyBit.scala 36:32]
  assign _GEN_134 = _GEN_791 | _GEN_110; // @[BusyBit.scala 36:32]
  assign _GEN_135 = _GEN_792 | _GEN_111; // @[BusyBit.scala 36:32]
  assign _GEN_137 = _T_31 ? _GEN_129 : _GEN_105; // @[BusyBit.scala 35:57]
  assign _GEN_138 = _T_31 ? _GEN_130 : _GEN_106; // @[BusyBit.scala 35:57]
  assign _GEN_139 = _T_31 ? _GEN_131 : _GEN_107; // @[BusyBit.scala 35:57]
  assign _GEN_140 = _T_31 ? _GEN_132 : _GEN_108; // @[BusyBit.scala 35:57]
  assign _GEN_141 = _T_31 ? _GEN_133 : _GEN_109; // @[BusyBit.scala 35:57]
  assign _GEN_142 = _T_31 ? _GEN_134 : _GEN_110; // @[BusyBit.scala 35:57]
  assign _GEN_143 = _T_31 ? _GEN_135 : _GEN_111; // @[BusyBit.scala 35:57]
  assign _GEN_145 = _T_29 ? _GEN_113 : _GEN_137; // @[BusyBit.scala 33:71]
  assign _GEN_146 = _T_29 ? _GEN_114 : _GEN_138; // @[BusyBit.scala 33:71]
  assign _GEN_147 = _T_29 ? _GEN_115 : _GEN_139; // @[BusyBit.scala 33:71]
  assign _GEN_148 = _T_29 ? _GEN_116 : _GEN_140; // @[BusyBit.scala 33:71]
  assign _GEN_149 = _T_29 ? _GEN_117 : _GEN_141; // @[BusyBit.scala 33:71]
  assign _GEN_150 = _T_29 ? _GEN_118 : _GEN_142; // @[BusyBit.scala 33:71]
  assign _GEN_151 = _T_29 ? _GEN_119 : _GEN_143; // @[BusyBit.scala 33:71]
  assign _GEN_153 = _T_17 ? _GEN_113 : _GEN_145; // @[BusyBit.scala 31:57]
  assign _GEN_154 = _T_17 ? _GEN_114 : _GEN_146; // @[BusyBit.scala 31:57]
  assign _GEN_155 = _T_17 ? _GEN_115 : _GEN_147; // @[BusyBit.scala 31:57]
  assign _GEN_156 = _T_17 ? _GEN_116 : _GEN_148; // @[BusyBit.scala 31:57]
  assign _GEN_157 = _T_17 ? _GEN_117 : _GEN_149; // @[BusyBit.scala 31:57]
  assign _GEN_158 = _T_17 ? _GEN_118 : _GEN_150; // @[BusyBit.scala 31:57]
  assign _GEN_159 = _T_17 ? _GEN_119 : _GEN_151; // @[BusyBit.scala 31:57]
  assign _GEN_161 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_153; // @[BusyBit.scala 32:39]
  assign _GEN_162 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_154; // @[BusyBit.scala 32:39]
  assign _GEN_163 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_155; // @[BusyBit.scala 32:39]
  assign _GEN_164 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_156; // @[BusyBit.scala 32:39]
  assign _GEN_165 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_157; // @[BusyBit.scala 32:39]
  assign _GEN_166 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_158; // @[BusyBit.scala 32:39]
  assign _GEN_167 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_159; // @[BusyBit.scala 32:39]
  assign _T_33 = io_release_0_rd_addr == 3'h3; // @[BusyBit.scala 33:62]
  assign _T_34 = io_release_0_rf_w & _T_33; // @[BusyBit.scala 33:37]
  assign _T_35 = io_req_rd_addr == 3'h3; // @[BusyBit.scala 35:48]
  assign _T_36 = io_req_rd_w & _T_35; // @[BusyBit.scala 35:30]
  assign _GEN_177 = _GEN_786 | _GEN_153; // @[BusyBit.scala 36:32]
  assign _GEN_178 = _GEN_787 | _GEN_154; // @[BusyBit.scala 36:32]
  assign _GEN_179 = _GEN_788 | _GEN_155; // @[BusyBit.scala 36:32]
  assign _GEN_180 = _GEN_789 | _GEN_156; // @[BusyBit.scala 36:32]
  assign _GEN_181 = _GEN_790 | _GEN_157; // @[BusyBit.scala 36:32]
  assign _GEN_182 = _GEN_791 | _GEN_158; // @[BusyBit.scala 36:32]
  assign _GEN_183 = _GEN_792 | _GEN_159; // @[BusyBit.scala 36:32]
  assign _GEN_185 = _T_36 ? _GEN_177 : _GEN_153; // @[BusyBit.scala 35:57]
  assign _GEN_186 = _T_36 ? _GEN_178 : _GEN_154; // @[BusyBit.scala 35:57]
  assign _GEN_187 = _T_36 ? _GEN_179 : _GEN_155; // @[BusyBit.scala 35:57]
  assign _GEN_188 = _T_36 ? _GEN_180 : _GEN_156; // @[BusyBit.scala 35:57]
  assign _GEN_189 = _T_36 ? _GEN_181 : _GEN_157; // @[BusyBit.scala 35:57]
  assign _GEN_190 = _T_36 ? _GEN_182 : _GEN_158; // @[BusyBit.scala 35:57]
  assign _GEN_191 = _T_36 ? _GEN_183 : _GEN_159; // @[BusyBit.scala 35:57]
  assign _GEN_193 = _T_34 ? _GEN_161 : _GEN_185; // @[BusyBit.scala 33:71]
  assign _GEN_194 = _T_34 ? _GEN_162 : _GEN_186; // @[BusyBit.scala 33:71]
  assign _GEN_195 = _T_34 ? _GEN_163 : _GEN_187; // @[BusyBit.scala 33:71]
  assign _GEN_196 = _T_34 ? _GEN_164 : _GEN_188; // @[BusyBit.scala 33:71]
  assign _GEN_197 = _T_34 ? _GEN_165 : _GEN_189; // @[BusyBit.scala 33:71]
  assign _GEN_198 = _T_34 ? _GEN_166 : _GEN_190; // @[BusyBit.scala 33:71]
  assign _GEN_199 = _T_34 ? _GEN_167 : _GEN_191; // @[BusyBit.scala 33:71]
  assign _GEN_201 = _T_17 ? _GEN_161 : _GEN_193; // @[BusyBit.scala 31:57]
  assign _GEN_202 = _T_17 ? _GEN_162 : _GEN_194; // @[BusyBit.scala 31:57]
  assign _GEN_203 = _T_17 ? _GEN_163 : _GEN_195; // @[BusyBit.scala 31:57]
  assign _GEN_204 = _T_17 ? _GEN_164 : _GEN_196; // @[BusyBit.scala 31:57]
  assign _GEN_205 = _T_17 ? _GEN_165 : _GEN_197; // @[BusyBit.scala 31:57]
  assign _GEN_206 = _T_17 ? _GEN_166 : _GEN_198; // @[BusyBit.scala 31:57]
  assign _GEN_207 = _T_17 ? _GEN_167 : _GEN_199; // @[BusyBit.scala 31:57]
  assign _GEN_209 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_201; // @[BusyBit.scala 32:39]
  assign _GEN_210 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_202; // @[BusyBit.scala 32:39]
  assign _GEN_211 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_203; // @[BusyBit.scala 32:39]
  assign _GEN_212 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_204; // @[BusyBit.scala 32:39]
  assign _GEN_213 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_205; // @[BusyBit.scala 32:39]
  assign _GEN_214 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_206; // @[BusyBit.scala 32:39]
  assign _GEN_215 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_207; // @[BusyBit.scala 32:39]
  assign _T_38 = io_release_0_rd_addr == 3'h4; // @[BusyBit.scala 33:62]
  assign _T_39 = io_release_0_rf_w & _T_38; // @[BusyBit.scala 33:37]
  assign _T_40 = io_req_rd_addr == 3'h4; // @[BusyBit.scala 35:48]
  assign _T_41 = io_req_rd_w & _T_40; // @[BusyBit.scala 35:30]
  assign _GEN_225 = _GEN_786 | _GEN_201; // @[BusyBit.scala 36:32]
  assign _GEN_226 = _GEN_787 | _GEN_202; // @[BusyBit.scala 36:32]
  assign _GEN_227 = _GEN_788 | _GEN_203; // @[BusyBit.scala 36:32]
  assign _GEN_228 = _GEN_789 | _GEN_204; // @[BusyBit.scala 36:32]
  assign _GEN_229 = _GEN_790 | _GEN_205; // @[BusyBit.scala 36:32]
  assign _GEN_230 = _GEN_791 | _GEN_206; // @[BusyBit.scala 36:32]
  assign _GEN_231 = _GEN_792 | _GEN_207; // @[BusyBit.scala 36:32]
  assign _GEN_233 = _T_41 ? _GEN_225 : _GEN_201; // @[BusyBit.scala 35:57]
  assign _GEN_234 = _T_41 ? _GEN_226 : _GEN_202; // @[BusyBit.scala 35:57]
  assign _GEN_235 = _T_41 ? _GEN_227 : _GEN_203; // @[BusyBit.scala 35:57]
  assign _GEN_236 = _T_41 ? _GEN_228 : _GEN_204; // @[BusyBit.scala 35:57]
  assign _GEN_237 = _T_41 ? _GEN_229 : _GEN_205; // @[BusyBit.scala 35:57]
  assign _GEN_238 = _T_41 ? _GEN_230 : _GEN_206; // @[BusyBit.scala 35:57]
  assign _GEN_239 = _T_41 ? _GEN_231 : _GEN_207; // @[BusyBit.scala 35:57]
  assign _GEN_241 = _T_39 ? _GEN_209 : _GEN_233; // @[BusyBit.scala 33:71]
  assign _GEN_242 = _T_39 ? _GEN_210 : _GEN_234; // @[BusyBit.scala 33:71]
  assign _GEN_243 = _T_39 ? _GEN_211 : _GEN_235; // @[BusyBit.scala 33:71]
  assign _GEN_244 = _T_39 ? _GEN_212 : _GEN_236; // @[BusyBit.scala 33:71]
  assign _GEN_245 = _T_39 ? _GEN_213 : _GEN_237; // @[BusyBit.scala 33:71]
  assign _GEN_246 = _T_39 ? _GEN_214 : _GEN_238; // @[BusyBit.scala 33:71]
  assign _GEN_247 = _T_39 ? _GEN_215 : _GEN_239; // @[BusyBit.scala 33:71]
  assign _GEN_249 = _T_17 ? _GEN_209 : _GEN_241; // @[BusyBit.scala 31:57]
  assign _GEN_250 = _T_17 ? _GEN_210 : _GEN_242; // @[BusyBit.scala 31:57]
  assign _GEN_251 = _T_17 ? _GEN_211 : _GEN_243; // @[BusyBit.scala 31:57]
  assign _GEN_252 = _T_17 ? _GEN_212 : _GEN_244; // @[BusyBit.scala 31:57]
  assign _GEN_253 = _T_17 ? _GEN_213 : _GEN_245; // @[BusyBit.scala 31:57]
  assign _GEN_254 = _T_17 ? _GEN_214 : _GEN_246; // @[BusyBit.scala 31:57]
  assign _GEN_255 = _T_17 ? _GEN_215 : _GEN_247; // @[BusyBit.scala 31:57]
  assign _GEN_257 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_249; // @[BusyBit.scala 32:39]
  assign _GEN_258 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_250; // @[BusyBit.scala 32:39]
  assign _GEN_259 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_251; // @[BusyBit.scala 32:39]
  assign _GEN_260 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_252; // @[BusyBit.scala 32:39]
  assign _GEN_261 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_253; // @[BusyBit.scala 32:39]
  assign _GEN_262 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_254; // @[BusyBit.scala 32:39]
  assign _GEN_263 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_255; // @[BusyBit.scala 32:39]
  assign _T_43 = io_release_0_rd_addr == 3'h5; // @[BusyBit.scala 33:62]
  assign _T_44 = io_release_0_rf_w & _T_43; // @[BusyBit.scala 33:37]
  assign _T_45 = io_req_rd_addr == 3'h5; // @[BusyBit.scala 35:48]
  assign _T_46 = io_req_rd_w & _T_45; // @[BusyBit.scala 35:30]
  assign _GEN_273 = _GEN_786 | _GEN_249; // @[BusyBit.scala 36:32]
  assign _GEN_274 = _GEN_787 | _GEN_250; // @[BusyBit.scala 36:32]
  assign _GEN_275 = _GEN_788 | _GEN_251; // @[BusyBit.scala 36:32]
  assign _GEN_276 = _GEN_789 | _GEN_252; // @[BusyBit.scala 36:32]
  assign _GEN_277 = _GEN_790 | _GEN_253; // @[BusyBit.scala 36:32]
  assign _GEN_278 = _GEN_791 | _GEN_254; // @[BusyBit.scala 36:32]
  assign _GEN_279 = _GEN_792 | _GEN_255; // @[BusyBit.scala 36:32]
  assign _GEN_281 = _T_46 ? _GEN_273 : _GEN_249; // @[BusyBit.scala 35:57]
  assign _GEN_282 = _T_46 ? _GEN_274 : _GEN_250; // @[BusyBit.scala 35:57]
  assign _GEN_283 = _T_46 ? _GEN_275 : _GEN_251; // @[BusyBit.scala 35:57]
  assign _GEN_284 = _T_46 ? _GEN_276 : _GEN_252; // @[BusyBit.scala 35:57]
  assign _GEN_285 = _T_46 ? _GEN_277 : _GEN_253; // @[BusyBit.scala 35:57]
  assign _GEN_286 = _T_46 ? _GEN_278 : _GEN_254; // @[BusyBit.scala 35:57]
  assign _GEN_287 = _T_46 ? _GEN_279 : _GEN_255; // @[BusyBit.scala 35:57]
  assign _GEN_289 = _T_44 ? _GEN_257 : _GEN_281; // @[BusyBit.scala 33:71]
  assign _GEN_290 = _T_44 ? _GEN_258 : _GEN_282; // @[BusyBit.scala 33:71]
  assign _GEN_291 = _T_44 ? _GEN_259 : _GEN_283; // @[BusyBit.scala 33:71]
  assign _GEN_292 = _T_44 ? _GEN_260 : _GEN_284; // @[BusyBit.scala 33:71]
  assign _GEN_293 = _T_44 ? _GEN_261 : _GEN_285; // @[BusyBit.scala 33:71]
  assign _GEN_294 = _T_44 ? _GEN_262 : _GEN_286; // @[BusyBit.scala 33:71]
  assign _GEN_295 = _T_44 ? _GEN_263 : _GEN_287; // @[BusyBit.scala 33:71]
  assign _GEN_297 = _T_17 ? _GEN_257 : _GEN_289; // @[BusyBit.scala 31:57]
  assign _GEN_298 = _T_17 ? _GEN_258 : _GEN_290; // @[BusyBit.scala 31:57]
  assign _GEN_299 = _T_17 ? _GEN_259 : _GEN_291; // @[BusyBit.scala 31:57]
  assign _GEN_300 = _T_17 ? _GEN_260 : _GEN_292; // @[BusyBit.scala 31:57]
  assign _GEN_301 = _T_17 ? _GEN_261 : _GEN_293; // @[BusyBit.scala 31:57]
  assign _GEN_302 = _T_17 ? _GEN_262 : _GEN_294; // @[BusyBit.scala 31:57]
  assign _GEN_303 = _T_17 ? _GEN_263 : _GEN_295; // @[BusyBit.scala 31:57]
  assign _GEN_305 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_297; // @[BusyBit.scala 32:39]
  assign _GEN_306 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_298; // @[BusyBit.scala 32:39]
  assign _GEN_307 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_299; // @[BusyBit.scala 32:39]
  assign _GEN_308 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_300; // @[BusyBit.scala 32:39]
  assign _GEN_309 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_301; // @[BusyBit.scala 32:39]
  assign _GEN_310 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_302; // @[BusyBit.scala 32:39]
  assign _GEN_311 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_303; // @[BusyBit.scala 32:39]
  assign _T_48 = io_release_0_rd_addr == 3'h6; // @[BusyBit.scala 33:62]
  assign _T_49 = io_release_0_rf_w & _T_48; // @[BusyBit.scala 33:37]
  assign _T_50 = io_req_rd_addr == 3'h6; // @[BusyBit.scala 35:48]
  assign _T_51 = io_req_rd_w & _T_50; // @[BusyBit.scala 35:30]
  assign _GEN_321 = _GEN_786 | _GEN_297; // @[BusyBit.scala 36:32]
  assign _GEN_322 = _GEN_787 | _GEN_298; // @[BusyBit.scala 36:32]
  assign _GEN_323 = _GEN_788 | _GEN_299; // @[BusyBit.scala 36:32]
  assign _GEN_324 = _GEN_789 | _GEN_300; // @[BusyBit.scala 36:32]
  assign _GEN_325 = _GEN_790 | _GEN_301; // @[BusyBit.scala 36:32]
  assign _GEN_326 = _GEN_791 | _GEN_302; // @[BusyBit.scala 36:32]
  assign _GEN_327 = _GEN_792 | _GEN_303; // @[BusyBit.scala 36:32]
  assign _GEN_329 = _T_51 ? _GEN_321 : _GEN_297; // @[BusyBit.scala 35:57]
  assign _GEN_330 = _T_51 ? _GEN_322 : _GEN_298; // @[BusyBit.scala 35:57]
  assign _GEN_331 = _T_51 ? _GEN_323 : _GEN_299; // @[BusyBit.scala 35:57]
  assign _GEN_332 = _T_51 ? _GEN_324 : _GEN_300; // @[BusyBit.scala 35:57]
  assign _GEN_333 = _T_51 ? _GEN_325 : _GEN_301; // @[BusyBit.scala 35:57]
  assign _GEN_334 = _T_51 ? _GEN_326 : _GEN_302; // @[BusyBit.scala 35:57]
  assign _GEN_335 = _T_51 ? _GEN_327 : _GEN_303; // @[BusyBit.scala 35:57]
  assign _GEN_337 = _T_49 ? _GEN_305 : _GEN_329; // @[BusyBit.scala 33:71]
  assign _GEN_338 = _T_49 ? _GEN_306 : _GEN_330; // @[BusyBit.scala 33:71]
  assign _GEN_339 = _T_49 ? _GEN_307 : _GEN_331; // @[BusyBit.scala 33:71]
  assign _GEN_340 = _T_49 ? _GEN_308 : _GEN_332; // @[BusyBit.scala 33:71]
  assign _GEN_341 = _T_49 ? _GEN_309 : _GEN_333; // @[BusyBit.scala 33:71]
  assign _GEN_342 = _T_49 ? _GEN_310 : _GEN_334; // @[BusyBit.scala 33:71]
  assign _GEN_343 = _T_49 ? _GEN_311 : _GEN_335; // @[BusyBit.scala 33:71]
  assign _GEN_345 = _T_17 ? _GEN_305 : _GEN_337; // @[BusyBit.scala 31:57]
  assign _GEN_346 = _T_17 ? _GEN_306 : _GEN_338; // @[BusyBit.scala 31:57]
  assign _GEN_347 = _T_17 ? _GEN_307 : _GEN_339; // @[BusyBit.scala 31:57]
  assign _GEN_348 = _T_17 ? _GEN_308 : _GEN_340; // @[BusyBit.scala 31:57]
  assign _GEN_349 = _T_17 ? _GEN_309 : _GEN_341; // @[BusyBit.scala 31:57]
  assign _GEN_350 = _T_17 ? _GEN_310 : _GEN_342; // @[BusyBit.scala 31:57]
  assign _GEN_351 = _T_17 ? _GEN_311 : _GEN_343; // @[BusyBit.scala 31:57]
  assign _GEN_353 = 3'h1 == io_release_0_rd_addr ? 1'h0 : _GEN_345; // @[BusyBit.scala 32:39]
  assign _GEN_354 = 3'h2 == io_release_0_rd_addr ? 1'h0 : _GEN_346; // @[BusyBit.scala 32:39]
  assign _GEN_355 = 3'h3 == io_release_0_rd_addr ? 1'h0 : _GEN_347; // @[BusyBit.scala 32:39]
  assign _GEN_356 = 3'h4 == io_release_0_rd_addr ? 1'h0 : _GEN_348; // @[BusyBit.scala 32:39]
  assign _GEN_357 = 3'h5 == io_release_0_rd_addr ? 1'h0 : _GEN_349; // @[BusyBit.scala 32:39]
  assign _GEN_358 = 3'h6 == io_release_0_rd_addr ? 1'h0 : _GEN_350; // @[BusyBit.scala 32:39]
  assign _GEN_359 = 3'h7 == io_release_0_rd_addr ? 1'h0 : _GEN_351; // @[BusyBit.scala 32:39]
  assign _T_53 = io_release_0_rd_addr == 3'h7; // @[BusyBit.scala 33:62]
  assign _T_54 = io_release_0_rf_w & _T_53; // @[BusyBit.scala 33:37]
  assign _T_55 = io_req_rd_addr == 3'h7; // @[BusyBit.scala 35:48]
  assign _T_56 = io_req_rd_w & _T_55; // @[BusyBit.scala 35:30]
  assign _GEN_369 = _GEN_786 | _GEN_345; // @[BusyBit.scala 36:32]
  assign _GEN_370 = _GEN_787 | _GEN_346; // @[BusyBit.scala 36:32]
  assign _GEN_371 = _GEN_788 | _GEN_347; // @[BusyBit.scala 36:32]
  assign _GEN_372 = _GEN_789 | _GEN_348; // @[BusyBit.scala 36:32]
  assign _GEN_373 = _GEN_790 | _GEN_349; // @[BusyBit.scala 36:32]
  assign _GEN_374 = _GEN_791 | _GEN_350; // @[BusyBit.scala 36:32]
  assign _GEN_375 = _GEN_792 | _GEN_351; // @[BusyBit.scala 36:32]
  assign _GEN_377 = _T_56 ? _GEN_369 : _GEN_345; // @[BusyBit.scala 35:57]
  assign _GEN_378 = _T_56 ? _GEN_370 : _GEN_346; // @[BusyBit.scala 35:57]
  assign _GEN_379 = _T_56 ? _GEN_371 : _GEN_347; // @[BusyBit.scala 35:57]
  assign _GEN_380 = _T_56 ? _GEN_372 : _GEN_348; // @[BusyBit.scala 35:57]
  assign _GEN_381 = _T_56 ? _GEN_373 : _GEN_349; // @[BusyBit.scala 35:57]
  assign _GEN_382 = _T_56 ? _GEN_374 : _GEN_350; // @[BusyBit.scala 35:57]
  assign _GEN_383 = _T_56 ? _GEN_375 : _GEN_351; // @[BusyBit.scala 35:57]
  assign _GEN_385 = _T_54 ? _GEN_353 : _GEN_377; // @[BusyBit.scala 33:71]
  assign _GEN_386 = _T_54 ? _GEN_354 : _GEN_378; // @[BusyBit.scala 33:71]
  assign _GEN_387 = _T_54 ? _GEN_355 : _GEN_379; // @[BusyBit.scala 33:71]
  assign _GEN_388 = _T_54 ? _GEN_356 : _GEN_380; // @[BusyBit.scala 33:71]
  assign _GEN_389 = _T_54 ? _GEN_357 : _GEN_381; // @[BusyBit.scala 33:71]
  assign _GEN_390 = _T_54 ? _GEN_358 : _GEN_382; // @[BusyBit.scala 33:71]
  assign _GEN_391 = _T_54 ? _GEN_359 : _GEN_383; // @[BusyBit.scala 33:71]
  assign _GEN_393 = _T_17 ? _GEN_353 : _GEN_385; // @[BusyBit.scala 31:57]
  assign _GEN_394 = _T_17 ? _GEN_354 : _GEN_386; // @[BusyBit.scala 31:57]
  assign _GEN_395 = _T_17 ? _GEN_355 : _GEN_387; // @[BusyBit.scala 31:57]
  assign _GEN_396 = _T_17 ? _GEN_356 : _GEN_388; // @[BusyBit.scala 31:57]
  assign _GEN_397 = _T_17 ? _GEN_357 : _GEN_389; // @[BusyBit.scala 31:57]
  assign _GEN_398 = _T_17 ? _GEN_358 : _GEN_390; // @[BusyBit.scala 31:57]
  assign _GEN_399 = _T_17 ? _GEN_359 : _GEN_391; // @[BusyBit.scala 31:57]
  assign _GEN_417 = _GEN_786 | _GEN_393; // @[BusyBit.scala 36:32]
  assign _GEN_418 = _GEN_787 | _GEN_394; // @[BusyBit.scala 36:32]
  assign _GEN_419 = _GEN_788 | _GEN_395; // @[BusyBit.scala 36:32]
  assign _GEN_420 = _GEN_789 | _GEN_396; // @[BusyBit.scala 36:32]
  assign _GEN_421 = _GEN_790 | _GEN_397; // @[BusyBit.scala 36:32]
  assign _GEN_422 = _GEN_791 | _GEN_398; // @[BusyBit.scala 36:32]
  assign _GEN_423 = _GEN_792 | _GEN_399; // @[BusyBit.scala 36:32]
  assign _GEN_425 = _T_21 ? _GEN_417 : _GEN_393; // @[BusyBit.scala 35:57]
  assign _GEN_426 = _T_21 ? _GEN_418 : _GEN_394; // @[BusyBit.scala 35:57]
  assign _GEN_427 = _T_21 ? _GEN_419 : _GEN_395; // @[BusyBit.scala 35:57]
  assign _GEN_428 = _T_21 ? _GEN_420 : _GEN_396; // @[BusyBit.scala 35:57]
  assign _GEN_429 = _T_21 ? _GEN_421 : _GEN_397; // @[BusyBit.scala 35:57]
  assign _GEN_430 = _T_21 ? _GEN_422 : _GEN_398; // @[BusyBit.scala 35:57]
  assign _GEN_431 = _T_21 ? _GEN_423 : _GEN_399; // @[BusyBit.scala 35:57]
  assign _GEN_441 = _T_17 ? _GEN_393 : _GEN_425; // @[BusyBit.scala 31:57]
  assign _GEN_442 = _T_17 ? _GEN_394 : _GEN_426; // @[BusyBit.scala 31:57]
  assign _GEN_443 = _T_17 ? _GEN_395 : _GEN_427; // @[BusyBit.scala 31:57]
  assign _GEN_444 = _T_17 ? _GEN_396 : _GEN_428; // @[BusyBit.scala 31:57]
  assign _GEN_445 = _T_17 ? _GEN_397 : _GEN_429; // @[BusyBit.scala 31:57]
  assign _GEN_446 = _T_17 ? _GEN_398 : _GEN_430; // @[BusyBit.scala 31:57]
  assign _GEN_447 = _T_17 ? _GEN_399 : _GEN_431; // @[BusyBit.scala 31:57]
  assign _GEN_465 = _GEN_786 | _GEN_441; // @[BusyBit.scala 36:32]
  assign _GEN_466 = _GEN_787 | _GEN_442; // @[BusyBit.scala 36:32]
  assign _GEN_467 = _GEN_788 | _GEN_443; // @[BusyBit.scala 36:32]
  assign _GEN_468 = _GEN_789 | _GEN_444; // @[BusyBit.scala 36:32]
  assign _GEN_469 = _GEN_790 | _GEN_445; // @[BusyBit.scala 36:32]
  assign _GEN_470 = _GEN_791 | _GEN_446; // @[BusyBit.scala 36:32]
  assign _GEN_471 = _GEN_792 | _GEN_447; // @[BusyBit.scala 36:32]
  assign _GEN_473 = _T_26 ? _GEN_465 : _GEN_441; // @[BusyBit.scala 35:57]
  assign _GEN_474 = _T_26 ? _GEN_466 : _GEN_442; // @[BusyBit.scala 35:57]
  assign _GEN_475 = _T_26 ? _GEN_467 : _GEN_443; // @[BusyBit.scala 35:57]
  assign _GEN_476 = _T_26 ? _GEN_468 : _GEN_444; // @[BusyBit.scala 35:57]
  assign _GEN_477 = _T_26 ? _GEN_469 : _GEN_445; // @[BusyBit.scala 35:57]
  assign _GEN_478 = _T_26 ? _GEN_470 : _GEN_446; // @[BusyBit.scala 35:57]
  assign _GEN_479 = _T_26 ? _GEN_471 : _GEN_447; // @[BusyBit.scala 35:57]
  assign _GEN_489 = _T_17 ? _GEN_441 : _GEN_473; // @[BusyBit.scala 31:57]
  assign _GEN_490 = _T_17 ? _GEN_442 : _GEN_474; // @[BusyBit.scala 31:57]
  assign _GEN_491 = _T_17 ? _GEN_443 : _GEN_475; // @[BusyBit.scala 31:57]
  assign _GEN_492 = _T_17 ? _GEN_444 : _GEN_476; // @[BusyBit.scala 31:57]
  assign _GEN_493 = _T_17 ? _GEN_445 : _GEN_477; // @[BusyBit.scala 31:57]
  assign _GEN_494 = _T_17 ? _GEN_446 : _GEN_478; // @[BusyBit.scala 31:57]
  assign _GEN_495 = _T_17 ? _GEN_447 : _GEN_479; // @[BusyBit.scala 31:57]
  assign _GEN_513 = _GEN_786 | _GEN_489; // @[BusyBit.scala 36:32]
  assign _GEN_514 = _GEN_787 | _GEN_490; // @[BusyBit.scala 36:32]
  assign _GEN_515 = _GEN_788 | _GEN_491; // @[BusyBit.scala 36:32]
  assign _GEN_516 = _GEN_789 | _GEN_492; // @[BusyBit.scala 36:32]
  assign _GEN_517 = _GEN_790 | _GEN_493; // @[BusyBit.scala 36:32]
  assign _GEN_518 = _GEN_791 | _GEN_494; // @[BusyBit.scala 36:32]
  assign _GEN_519 = _GEN_792 | _GEN_495; // @[BusyBit.scala 36:32]
  assign _GEN_521 = _T_31 ? _GEN_513 : _GEN_489; // @[BusyBit.scala 35:57]
  assign _GEN_522 = _T_31 ? _GEN_514 : _GEN_490; // @[BusyBit.scala 35:57]
  assign _GEN_523 = _T_31 ? _GEN_515 : _GEN_491; // @[BusyBit.scala 35:57]
  assign _GEN_524 = _T_31 ? _GEN_516 : _GEN_492; // @[BusyBit.scala 35:57]
  assign _GEN_525 = _T_31 ? _GEN_517 : _GEN_493; // @[BusyBit.scala 35:57]
  assign _GEN_526 = _T_31 ? _GEN_518 : _GEN_494; // @[BusyBit.scala 35:57]
  assign _GEN_527 = _T_31 ? _GEN_519 : _GEN_495; // @[BusyBit.scala 35:57]
  assign _GEN_537 = _T_17 ? _GEN_489 : _GEN_521; // @[BusyBit.scala 31:57]
  assign _GEN_538 = _T_17 ? _GEN_490 : _GEN_522; // @[BusyBit.scala 31:57]
  assign _GEN_539 = _T_17 ? _GEN_491 : _GEN_523; // @[BusyBit.scala 31:57]
  assign _GEN_540 = _T_17 ? _GEN_492 : _GEN_524; // @[BusyBit.scala 31:57]
  assign _GEN_541 = _T_17 ? _GEN_493 : _GEN_525; // @[BusyBit.scala 31:57]
  assign _GEN_542 = _T_17 ? _GEN_494 : _GEN_526; // @[BusyBit.scala 31:57]
  assign _GEN_543 = _T_17 ? _GEN_495 : _GEN_527; // @[BusyBit.scala 31:57]
  assign _GEN_561 = _GEN_786 | _GEN_537; // @[BusyBit.scala 36:32]
  assign _GEN_562 = _GEN_787 | _GEN_538; // @[BusyBit.scala 36:32]
  assign _GEN_563 = _GEN_788 | _GEN_539; // @[BusyBit.scala 36:32]
  assign _GEN_564 = _GEN_789 | _GEN_540; // @[BusyBit.scala 36:32]
  assign _GEN_565 = _GEN_790 | _GEN_541; // @[BusyBit.scala 36:32]
  assign _GEN_566 = _GEN_791 | _GEN_542; // @[BusyBit.scala 36:32]
  assign _GEN_567 = _GEN_792 | _GEN_543; // @[BusyBit.scala 36:32]
  assign _GEN_569 = _T_36 ? _GEN_561 : _GEN_537; // @[BusyBit.scala 35:57]
  assign _GEN_570 = _T_36 ? _GEN_562 : _GEN_538; // @[BusyBit.scala 35:57]
  assign _GEN_571 = _T_36 ? _GEN_563 : _GEN_539; // @[BusyBit.scala 35:57]
  assign _GEN_572 = _T_36 ? _GEN_564 : _GEN_540; // @[BusyBit.scala 35:57]
  assign _GEN_573 = _T_36 ? _GEN_565 : _GEN_541; // @[BusyBit.scala 35:57]
  assign _GEN_574 = _T_36 ? _GEN_566 : _GEN_542; // @[BusyBit.scala 35:57]
  assign _GEN_575 = _T_36 ? _GEN_567 : _GEN_543; // @[BusyBit.scala 35:57]
  assign _GEN_585 = _T_17 ? _GEN_537 : _GEN_569; // @[BusyBit.scala 31:57]
  assign _GEN_586 = _T_17 ? _GEN_538 : _GEN_570; // @[BusyBit.scala 31:57]
  assign _GEN_587 = _T_17 ? _GEN_539 : _GEN_571; // @[BusyBit.scala 31:57]
  assign _GEN_588 = _T_17 ? _GEN_540 : _GEN_572; // @[BusyBit.scala 31:57]
  assign _GEN_589 = _T_17 ? _GEN_541 : _GEN_573; // @[BusyBit.scala 31:57]
  assign _GEN_590 = _T_17 ? _GEN_542 : _GEN_574; // @[BusyBit.scala 31:57]
  assign _GEN_591 = _T_17 ? _GEN_543 : _GEN_575; // @[BusyBit.scala 31:57]
  assign _GEN_609 = _GEN_786 | _GEN_585; // @[BusyBit.scala 36:32]
  assign _GEN_610 = _GEN_787 | _GEN_586; // @[BusyBit.scala 36:32]
  assign _GEN_611 = _GEN_788 | _GEN_587; // @[BusyBit.scala 36:32]
  assign _GEN_612 = _GEN_789 | _GEN_588; // @[BusyBit.scala 36:32]
  assign _GEN_613 = _GEN_790 | _GEN_589; // @[BusyBit.scala 36:32]
  assign _GEN_614 = _GEN_791 | _GEN_590; // @[BusyBit.scala 36:32]
  assign _GEN_615 = _GEN_792 | _GEN_591; // @[BusyBit.scala 36:32]
  assign _GEN_617 = _T_41 ? _GEN_609 : _GEN_585; // @[BusyBit.scala 35:57]
  assign _GEN_618 = _T_41 ? _GEN_610 : _GEN_586; // @[BusyBit.scala 35:57]
  assign _GEN_619 = _T_41 ? _GEN_611 : _GEN_587; // @[BusyBit.scala 35:57]
  assign _GEN_620 = _T_41 ? _GEN_612 : _GEN_588; // @[BusyBit.scala 35:57]
  assign _GEN_621 = _T_41 ? _GEN_613 : _GEN_589; // @[BusyBit.scala 35:57]
  assign _GEN_622 = _T_41 ? _GEN_614 : _GEN_590; // @[BusyBit.scala 35:57]
  assign _GEN_623 = _T_41 ? _GEN_615 : _GEN_591; // @[BusyBit.scala 35:57]
  assign _GEN_633 = _T_17 ? _GEN_585 : _GEN_617; // @[BusyBit.scala 31:57]
  assign _GEN_634 = _T_17 ? _GEN_586 : _GEN_618; // @[BusyBit.scala 31:57]
  assign _GEN_635 = _T_17 ? _GEN_587 : _GEN_619; // @[BusyBit.scala 31:57]
  assign _GEN_636 = _T_17 ? _GEN_588 : _GEN_620; // @[BusyBit.scala 31:57]
  assign _GEN_637 = _T_17 ? _GEN_589 : _GEN_621; // @[BusyBit.scala 31:57]
  assign _GEN_638 = _T_17 ? _GEN_590 : _GEN_622; // @[BusyBit.scala 31:57]
  assign _GEN_639 = _T_17 ? _GEN_591 : _GEN_623; // @[BusyBit.scala 31:57]
  assign _GEN_657 = _GEN_786 | _GEN_633; // @[BusyBit.scala 36:32]
  assign _GEN_658 = _GEN_787 | _GEN_634; // @[BusyBit.scala 36:32]
  assign _GEN_659 = _GEN_788 | _GEN_635; // @[BusyBit.scala 36:32]
  assign _GEN_660 = _GEN_789 | _GEN_636; // @[BusyBit.scala 36:32]
  assign _GEN_661 = _GEN_790 | _GEN_637; // @[BusyBit.scala 36:32]
  assign _GEN_662 = _GEN_791 | _GEN_638; // @[BusyBit.scala 36:32]
  assign _GEN_663 = _GEN_792 | _GEN_639; // @[BusyBit.scala 36:32]
  assign _GEN_665 = _T_46 ? _GEN_657 : _GEN_633; // @[BusyBit.scala 35:57]
  assign _GEN_666 = _T_46 ? _GEN_658 : _GEN_634; // @[BusyBit.scala 35:57]
  assign _GEN_667 = _T_46 ? _GEN_659 : _GEN_635; // @[BusyBit.scala 35:57]
  assign _GEN_668 = _T_46 ? _GEN_660 : _GEN_636; // @[BusyBit.scala 35:57]
  assign _GEN_669 = _T_46 ? _GEN_661 : _GEN_637; // @[BusyBit.scala 35:57]
  assign _GEN_670 = _T_46 ? _GEN_662 : _GEN_638; // @[BusyBit.scala 35:57]
  assign _GEN_671 = _T_46 ? _GEN_663 : _GEN_639; // @[BusyBit.scala 35:57]
  assign _GEN_681 = _T_17 ? _GEN_633 : _GEN_665; // @[BusyBit.scala 31:57]
  assign _GEN_682 = _T_17 ? _GEN_634 : _GEN_666; // @[BusyBit.scala 31:57]
  assign _GEN_683 = _T_17 ? _GEN_635 : _GEN_667; // @[BusyBit.scala 31:57]
  assign _GEN_684 = _T_17 ? _GEN_636 : _GEN_668; // @[BusyBit.scala 31:57]
  assign _GEN_685 = _T_17 ? _GEN_637 : _GEN_669; // @[BusyBit.scala 31:57]
  assign _GEN_686 = _T_17 ? _GEN_638 : _GEN_670; // @[BusyBit.scala 31:57]
  assign _GEN_687 = _T_17 ? _GEN_639 : _GEN_671; // @[BusyBit.scala 31:57]
  assign _GEN_705 = _GEN_786 | _GEN_681; // @[BusyBit.scala 36:32]
  assign _GEN_706 = _GEN_787 | _GEN_682; // @[BusyBit.scala 36:32]
  assign _GEN_707 = _GEN_788 | _GEN_683; // @[BusyBit.scala 36:32]
  assign _GEN_708 = _GEN_789 | _GEN_684; // @[BusyBit.scala 36:32]
  assign _GEN_709 = _GEN_790 | _GEN_685; // @[BusyBit.scala 36:32]
  assign _GEN_710 = _GEN_791 | _GEN_686; // @[BusyBit.scala 36:32]
  assign _GEN_711 = _GEN_792 | _GEN_687; // @[BusyBit.scala 36:32]
  assign _GEN_713 = _T_51 ? _GEN_705 : _GEN_681; // @[BusyBit.scala 35:57]
  assign _GEN_714 = _T_51 ? _GEN_706 : _GEN_682; // @[BusyBit.scala 35:57]
  assign _GEN_715 = _T_51 ? _GEN_707 : _GEN_683; // @[BusyBit.scala 35:57]
  assign _GEN_716 = _T_51 ? _GEN_708 : _GEN_684; // @[BusyBit.scala 35:57]
  assign _GEN_717 = _T_51 ? _GEN_709 : _GEN_685; // @[BusyBit.scala 35:57]
  assign _GEN_718 = _T_51 ? _GEN_710 : _GEN_686; // @[BusyBit.scala 35:57]
  assign _GEN_719 = _T_51 ? _GEN_711 : _GEN_687; // @[BusyBit.scala 35:57]
  assign _GEN_729 = _T_17 ? _GEN_681 : _GEN_713; // @[BusyBit.scala 31:57]
  assign _GEN_730 = _T_17 ? _GEN_682 : _GEN_714; // @[BusyBit.scala 31:57]
  assign _GEN_731 = _T_17 ? _GEN_683 : _GEN_715; // @[BusyBit.scala 31:57]
  assign _GEN_732 = _T_17 ? _GEN_684 : _GEN_716; // @[BusyBit.scala 31:57]
  assign _GEN_733 = _T_17 ? _GEN_685 : _GEN_717; // @[BusyBit.scala 31:57]
  assign _GEN_734 = _T_17 ? _GEN_686 : _GEN_718; // @[BusyBit.scala 31:57]
  assign _GEN_735 = _T_17 ? _GEN_687 : _GEN_719; // @[BusyBit.scala 31:57]
  assign _GEN_753 = _GEN_786 | _GEN_729; // @[BusyBit.scala 36:32]
  assign _GEN_754 = _GEN_787 | _GEN_730; // @[BusyBit.scala 36:32]
  assign _GEN_755 = _GEN_788 | _GEN_731; // @[BusyBit.scala 36:32]
  assign _GEN_756 = _GEN_789 | _GEN_732; // @[BusyBit.scala 36:32]
  assign _GEN_757 = _GEN_790 | _GEN_733; // @[BusyBit.scala 36:32]
  assign _GEN_758 = _GEN_791 | _GEN_734; // @[BusyBit.scala 36:32]
  assign _GEN_759 = _GEN_792 | _GEN_735; // @[BusyBit.scala 36:32]
  assign _T_97 = $unsigned(reset); // @[BusyBit.scala 40:9]
  assign _T_98 = _T_97 == 1'h0; // @[BusyBit.scala 40:9]
  assign io_rs_available_0 = _T_7 | _T_2; // @[BusyBit.scala 27:24]
  assign io_rs_available_1 = _T_15 | _T_10; // @[BusyBit.scala 27:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy_bit_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  busy_bit_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  busy_bit_3 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  busy_bit_4 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  busy_bit_5 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  busy_bit_6 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  busy_bit_7 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      busy_bit_1 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h1 == io_release_0_rd_addr) begin
                        busy_bit_1 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h1 == io_release_0_rd_addr) begin
                          busy_bit_1 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h1 == io_release_0_rd_addr) begin
                            busy_bit_1 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h1 == io_release_0_rd_addr) begin
                              busy_bit_1 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h1 == io_release_0_rd_addr) begin
                                busy_bit_1 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h1 == io_release_0_rd_addr) begin
                                  busy_bit_1 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h1 == io_release_0_rd_addr) begin
                                    busy_bit_1 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h1 == io_release_0_rd_addr) begin
                                      busy_bit_1 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h1 == io_release_0_rd_addr) begin
                                      busy_bit_1 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_1 <= _GEN_33;
                                  end
                                end else if (_T_24) begin
                                  if (3'h1 == io_release_0_rd_addr) begin
                                    busy_bit_1 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h1 == io_release_0_rd_addr) begin
                                      busy_bit_1 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h1 == io_release_0_rd_addr) begin
                                      busy_bit_1 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_1 <= _GEN_33;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_1 <= _GEN_81;
                                end else if (_T_17) begin
                                  busy_bit_1 <= _GEN_17;
                                end else if (_T_19) begin
                                  busy_bit_1 <= _GEN_17;
                                end else if (_T_21) begin
                                  busy_bit_1 <= _GEN_33;
                                end
                              end else if (_T_29) begin
                                if (3'h1 == io_release_0_rd_addr) begin
                                  busy_bit_1 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h1 == io_release_0_rd_addr) begin
                                    busy_bit_1 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_1 <= _GEN_17;
                                  end else if (_T_19) begin
                                    busy_bit_1 <= _GEN_17;
                                  end else if (_T_21) begin
                                    busy_bit_1 <= _GEN_33;
                                  end
                                end else if (_T_24) begin
                                  if (3'h1 == io_release_0_rd_addr) begin
                                    busy_bit_1 <= 1'h0;
                                  end else begin
                                    busy_bit_1 <= _GEN_57;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_1 <= _GEN_81;
                                end else begin
                                  busy_bit_1 <= _GEN_57;
                                end
                              end else if (_T_31) begin
                                busy_bit_1 <= _GEN_129;
                              end else if (_T_17) begin
                                busy_bit_1 <= _GEN_65;
                              end else if (_T_24) begin
                                busy_bit_1 <= _GEN_65;
                              end else if (_T_26) begin
                                busy_bit_1 <= _GEN_81;
                              end else begin
                                busy_bit_1 <= _GEN_57;
                              end
                            end else if (_T_34) begin
                              if (3'h1 == io_release_0_rd_addr) begin
                                busy_bit_1 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h1 == io_release_0_rd_addr) begin
                                  busy_bit_1 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_1 <= _GEN_65;
                                end else if (_T_24) begin
                                  busy_bit_1 <= _GEN_65;
                                end else if (_T_26) begin
                                  busy_bit_1 <= _GEN_81;
                                end else begin
                                  busy_bit_1 <= _GEN_57;
                                end
                              end else if (_T_29) begin
                                if (3'h1 == io_release_0_rd_addr) begin
                                  busy_bit_1 <= 1'h0;
                                end else begin
                                  busy_bit_1 <= _GEN_105;
                                end
                              end else if (_T_31) begin
                                busy_bit_1 <= _GEN_129;
                              end else begin
                                busy_bit_1 <= _GEN_105;
                              end
                            end else if (_T_36) begin
                              busy_bit_1 <= _GEN_177;
                            end else if (_T_17) begin
                              busy_bit_1 <= _GEN_113;
                            end else if (_T_29) begin
                              busy_bit_1 <= _GEN_113;
                            end else if (_T_31) begin
                              busy_bit_1 <= _GEN_129;
                            end else begin
                              busy_bit_1 <= _GEN_105;
                            end
                          end else if (_T_39) begin
                            if (3'h1 == io_release_0_rd_addr) begin
                              busy_bit_1 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h1 == io_release_0_rd_addr) begin
                                busy_bit_1 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_1 <= _GEN_113;
                              end else if (_T_29) begin
                                busy_bit_1 <= _GEN_113;
                              end else if (_T_31) begin
                                busy_bit_1 <= _GEN_129;
                              end else begin
                                busy_bit_1 <= _GEN_105;
                              end
                            end else if (_T_34) begin
                              if (3'h1 == io_release_0_rd_addr) begin
                                busy_bit_1 <= 1'h0;
                              end else begin
                                busy_bit_1 <= _GEN_153;
                              end
                            end else if (_T_36) begin
                              busy_bit_1 <= _GEN_177;
                            end else begin
                              busy_bit_1 <= _GEN_153;
                            end
                          end else if (_T_41) begin
                            busy_bit_1 <= _GEN_225;
                          end else if (_T_17) begin
                            busy_bit_1 <= _GEN_161;
                          end else if (_T_34) begin
                            busy_bit_1 <= _GEN_161;
                          end else if (_T_36) begin
                            busy_bit_1 <= _GEN_177;
                          end else begin
                            busy_bit_1 <= _GEN_153;
                          end
                        end else if (_T_44) begin
                          if (3'h1 == io_release_0_rd_addr) begin
                            busy_bit_1 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h1 == io_release_0_rd_addr) begin
                              busy_bit_1 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_1 <= _GEN_161;
                            end else if (_T_34) begin
                              busy_bit_1 <= _GEN_161;
                            end else if (_T_36) begin
                              busy_bit_1 <= _GEN_177;
                            end else begin
                              busy_bit_1 <= _GEN_153;
                            end
                          end else if (_T_39) begin
                            if (3'h1 == io_release_0_rd_addr) begin
                              busy_bit_1 <= 1'h0;
                            end else begin
                              busy_bit_1 <= _GEN_201;
                            end
                          end else if (_T_41) begin
                            busy_bit_1 <= _GEN_225;
                          end else begin
                            busy_bit_1 <= _GEN_201;
                          end
                        end else if (_T_46) begin
                          busy_bit_1 <= _GEN_273;
                        end else if (_T_17) begin
                          busy_bit_1 <= _GEN_209;
                        end else if (_T_39) begin
                          busy_bit_1 <= _GEN_209;
                        end else if (_T_41) begin
                          busy_bit_1 <= _GEN_225;
                        end else begin
                          busy_bit_1 <= _GEN_201;
                        end
                      end else if (_T_49) begin
                        if (3'h1 == io_release_0_rd_addr) begin
                          busy_bit_1 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h1 == io_release_0_rd_addr) begin
                            busy_bit_1 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_1 <= _GEN_209;
                          end else if (_T_39) begin
                            busy_bit_1 <= _GEN_209;
                          end else if (_T_41) begin
                            busy_bit_1 <= _GEN_225;
                          end else begin
                            busy_bit_1 <= _GEN_201;
                          end
                        end else if (_T_44) begin
                          if (3'h1 == io_release_0_rd_addr) begin
                            busy_bit_1 <= 1'h0;
                          end else begin
                            busy_bit_1 <= _GEN_249;
                          end
                        end else if (_T_46) begin
                          busy_bit_1 <= _GEN_273;
                        end else begin
                          busy_bit_1 <= _GEN_249;
                        end
                      end else if (_T_51) begin
                        busy_bit_1 <= _GEN_321;
                      end else if (_T_17) begin
                        busy_bit_1 <= _GEN_257;
                      end else if (_T_44) begin
                        busy_bit_1 <= _GEN_257;
                      end else if (_T_46) begin
                        busy_bit_1 <= _GEN_273;
                      end else begin
                        busy_bit_1 <= _GEN_249;
                      end
                    end else if (_T_54) begin
                      if (3'h1 == io_release_0_rd_addr) begin
                        busy_bit_1 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h1 == io_release_0_rd_addr) begin
                          busy_bit_1 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_1 <= _GEN_257;
                        end else if (_T_44) begin
                          busy_bit_1 <= _GEN_257;
                        end else if (_T_46) begin
                          busy_bit_1 <= _GEN_273;
                        end else begin
                          busy_bit_1 <= _GEN_249;
                        end
                      end else if (_T_49) begin
                        if (3'h1 == io_release_0_rd_addr) begin
                          busy_bit_1 <= 1'h0;
                        end else begin
                          busy_bit_1 <= _GEN_297;
                        end
                      end else if (_T_51) begin
                        busy_bit_1 <= _GEN_321;
                      end else begin
                        busy_bit_1 <= _GEN_297;
                      end
                    end else if (_T_56) begin
                      busy_bit_1 <= _GEN_369;
                    end else if (_T_17) begin
                      busy_bit_1 <= _GEN_305;
                    end else if (_T_49) begin
                      busy_bit_1 <= _GEN_305;
                    end else if (_T_51) begin
                      busy_bit_1 <= _GEN_321;
                    end else begin
                      busy_bit_1 <= _GEN_297;
                    end
                  end else if (_T_21) begin
                    busy_bit_1 <= _GEN_417;
                  end else if (_T_17) begin
                    if (3'h1 == io_release_0_rd_addr) begin
                      busy_bit_1 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_1 <= _GEN_305;
                    end else if (_T_49) begin
                      busy_bit_1 <= _GEN_305;
                    end else if (_T_51) begin
                      busy_bit_1 <= _GEN_321;
                    end else begin
                      busy_bit_1 <= _GEN_297;
                    end
                  end else if (_T_54) begin
                    if (3'h1 == io_release_0_rd_addr) begin
                      busy_bit_1 <= 1'h0;
                    end else begin
                      busy_bit_1 <= _GEN_345;
                    end
                  end else if (_T_56) begin
                    busy_bit_1 <= _GEN_369;
                  end else begin
                    busy_bit_1 <= _GEN_345;
                  end
                end else if (_T_26) begin
                  busy_bit_1 <= _GEN_465;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_1 <= _GEN_353;
                  end else if (_T_54) begin
                    busy_bit_1 <= _GEN_353;
                  end else if (_T_56) begin
                    busy_bit_1 <= _GEN_369;
                  end else begin
                    busy_bit_1 <= _GEN_345;
                  end
                end else if (_T_21) begin
                  busy_bit_1 <= _GEN_417;
                end else if (_T_17) begin
                  busy_bit_1 <= _GEN_353;
                end else if (_T_54) begin
                  busy_bit_1 <= _GEN_353;
                end else if (_T_56) begin
                  busy_bit_1 <= _GEN_369;
                end else begin
                  busy_bit_1 <= _GEN_345;
                end
              end else if (_T_31) begin
                busy_bit_1 <= _GEN_513;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_1 <= _GEN_393;
                end else if (_T_21) begin
                  busy_bit_1 <= _GEN_417;
                end else begin
                  busy_bit_1 <= _GEN_393;
                end
              end else if (_T_26) begin
                busy_bit_1 <= _GEN_465;
              end else if (_T_17) begin
                busy_bit_1 <= _GEN_393;
              end else if (_T_21) begin
                busy_bit_1 <= _GEN_417;
              end else begin
                busy_bit_1 <= _GEN_393;
              end
            end else if (_T_36) begin
              busy_bit_1 <= _GEN_561;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_1 <= _GEN_441;
              end else if (_T_26) begin
                busy_bit_1 <= _GEN_465;
              end else begin
                busy_bit_1 <= _GEN_441;
              end
            end else if (_T_31) begin
              busy_bit_1 <= _GEN_513;
            end else if (_T_17) begin
              busy_bit_1 <= _GEN_441;
            end else if (_T_26) begin
              busy_bit_1 <= _GEN_465;
            end else begin
              busy_bit_1 <= _GEN_441;
            end
          end else if (_T_41) begin
            busy_bit_1 <= _GEN_609;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_1 <= _GEN_489;
            end else if (_T_31) begin
              busy_bit_1 <= _GEN_513;
            end else begin
              busy_bit_1 <= _GEN_489;
            end
          end else if (_T_36) begin
            busy_bit_1 <= _GEN_561;
          end else if (_T_17) begin
            busy_bit_1 <= _GEN_489;
          end else if (_T_31) begin
            busy_bit_1 <= _GEN_513;
          end else begin
            busy_bit_1 <= _GEN_489;
          end
        end else if (_T_46) begin
          busy_bit_1 <= _GEN_657;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_1 <= _GEN_537;
          end else if (_T_36) begin
            busy_bit_1 <= _GEN_561;
          end else begin
            busy_bit_1 <= _GEN_537;
          end
        end else if (_T_41) begin
          busy_bit_1 <= _GEN_609;
        end else if (_T_17) begin
          busy_bit_1 <= _GEN_537;
        end else if (_T_36) begin
          busy_bit_1 <= _GEN_561;
        end else begin
          busy_bit_1 <= _GEN_537;
        end
      end else if (_T_51) begin
        busy_bit_1 <= _GEN_705;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_1 <= _GEN_585;
        end else if (_T_41) begin
          busy_bit_1 <= _GEN_609;
        end else begin
          busy_bit_1 <= _GEN_585;
        end
      end else if (_T_46) begin
        busy_bit_1 <= _GEN_657;
      end else if (_T_17) begin
        busy_bit_1 <= _GEN_585;
      end else if (_T_41) begin
        busy_bit_1 <= _GEN_609;
      end else begin
        busy_bit_1 <= _GEN_585;
      end
    end else if (_T_56) begin
      busy_bit_1 <= _GEN_753;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_1 <= _GEN_633;
      end else if (_T_46) begin
        busy_bit_1 <= _GEN_657;
      end else begin
        busy_bit_1 <= _GEN_633;
      end
    end else if (_T_51) begin
      busy_bit_1 <= _GEN_705;
    end else if (_T_17) begin
      busy_bit_1 <= _GEN_633;
    end else if (_T_46) begin
      busy_bit_1 <= _GEN_657;
    end else begin
      busy_bit_1 <= _GEN_633;
    end
    if (reset) begin
      busy_bit_2 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h2 == io_release_0_rd_addr) begin
                        busy_bit_2 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h2 == io_release_0_rd_addr) begin
                          busy_bit_2 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h2 == io_release_0_rd_addr) begin
                            busy_bit_2 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h2 == io_release_0_rd_addr) begin
                              busy_bit_2 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h2 == io_release_0_rd_addr) begin
                                busy_bit_2 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h2 == io_release_0_rd_addr) begin
                                  busy_bit_2 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h2 == io_release_0_rd_addr) begin
                                    busy_bit_2 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h2 == io_release_0_rd_addr) begin
                                      busy_bit_2 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h2 == io_release_0_rd_addr) begin
                                      busy_bit_2 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_2 <= _GEN_34;
                                  end
                                end else if (_T_24) begin
                                  if (3'h2 == io_release_0_rd_addr) begin
                                    busy_bit_2 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h2 == io_release_0_rd_addr) begin
                                      busy_bit_2 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h2 == io_release_0_rd_addr) begin
                                      busy_bit_2 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_2 <= _GEN_34;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_2 <= _GEN_82;
                                end else if (_T_17) begin
                                  busy_bit_2 <= _GEN_18;
                                end else if (_T_19) begin
                                  busy_bit_2 <= _GEN_18;
                                end else if (_T_21) begin
                                  busy_bit_2 <= _GEN_34;
                                end
                              end else if (_T_29) begin
                                if (3'h2 == io_release_0_rd_addr) begin
                                  busy_bit_2 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h2 == io_release_0_rd_addr) begin
                                    busy_bit_2 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_2 <= _GEN_18;
                                  end else if (_T_19) begin
                                    busy_bit_2 <= _GEN_18;
                                  end else if (_T_21) begin
                                    busy_bit_2 <= _GEN_34;
                                  end
                                end else if (_T_24) begin
                                  if (3'h2 == io_release_0_rd_addr) begin
                                    busy_bit_2 <= 1'h0;
                                  end else begin
                                    busy_bit_2 <= _GEN_58;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_2 <= _GEN_82;
                                end else begin
                                  busy_bit_2 <= _GEN_58;
                                end
                              end else if (_T_31) begin
                                busy_bit_2 <= _GEN_130;
                              end else if (_T_17) begin
                                busy_bit_2 <= _GEN_66;
                              end else if (_T_24) begin
                                busy_bit_2 <= _GEN_66;
                              end else if (_T_26) begin
                                busy_bit_2 <= _GEN_82;
                              end else begin
                                busy_bit_2 <= _GEN_58;
                              end
                            end else if (_T_34) begin
                              if (3'h2 == io_release_0_rd_addr) begin
                                busy_bit_2 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h2 == io_release_0_rd_addr) begin
                                  busy_bit_2 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_2 <= _GEN_66;
                                end else if (_T_24) begin
                                  busy_bit_2 <= _GEN_66;
                                end else if (_T_26) begin
                                  busy_bit_2 <= _GEN_82;
                                end else begin
                                  busy_bit_2 <= _GEN_58;
                                end
                              end else if (_T_29) begin
                                if (3'h2 == io_release_0_rd_addr) begin
                                  busy_bit_2 <= 1'h0;
                                end else begin
                                  busy_bit_2 <= _GEN_106;
                                end
                              end else if (_T_31) begin
                                busy_bit_2 <= _GEN_130;
                              end else begin
                                busy_bit_2 <= _GEN_106;
                              end
                            end else if (_T_36) begin
                              busy_bit_2 <= _GEN_178;
                            end else if (_T_17) begin
                              busy_bit_2 <= _GEN_114;
                            end else if (_T_29) begin
                              busy_bit_2 <= _GEN_114;
                            end else if (_T_31) begin
                              busy_bit_2 <= _GEN_130;
                            end else begin
                              busy_bit_2 <= _GEN_106;
                            end
                          end else if (_T_39) begin
                            if (3'h2 == io_release_0_rd_addr) begin
                              busy_bit_2 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h2 == io_release_0_rd_addr) begin
                                busy_bit_2 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_2 <= _GEN_114;
                              end else if (_T_29) begin
                                busy_bit_2 <= _GEN_114;
                              end else if (_T_31) begin
                                busy_bit_2 <= _GEN_130;
                              end else begin
                                busy_bit_2 <= _GEN_106;
                              end
                            end else if (_T_34) begin
                              if (3'h2 == io_release_0_rd_addr) begin
                                busy_bit_2 <= 1'h0;
                              end else begin
                                busy_bit_2 <= _GEN_154;
                              end
                            end else if (_T_36) begin
                              busy_bit_2 <= _GEN_178;
                            end else begin
                              busy_bit_2 <= _GEN_154;
                            end
                          end else if (_T_41) begin
                            busy_bit_2 <= _GEN_226;
                          end else if (_T_17) begin
                            busy_bit_2 <= _GEN_162;
                          end else if (_T_34) begin
                            busy_bit_2 <= _GEN_162;
                          end else if (_T_36) begin
                            busy_bit_2 <= _GEN_178;
                          end else begin
                            busy_bit_2 <= _GEN_154;
                          end
                        end else if (_T_44) begin
                          if (3'h2 == io_release_0_rd_addr) begin
                            busy_bit_2 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h2 == io_release_0_rd_addr) begin
                              busy_bit_2 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_2 <= _GEN_162;
                            end else if (_T_34) begin
                              busy_bit_2 <= _GEN_162;
                            end else if (_T_36) begin
                              busy_bit_2 <= _GEN_178;
                            end else begin
                              busy_bit_2 <= _GEN_154;
                            end
                          end else if (_T_39) begin
                            if (3'h2 == io_release_0_rd_addr) begin
                              busy_bit_2 <= 1'h0;
                            end else begin
                              busy_bit_2 <= _GEN_202;
                            end
                          end else if (_T_41) begin
                            busy_bit_2 <= _GEN_226;
                          end else begin
                            busy_bit_2 <= _GEN_202;
                          end
                        end else if (_T_46) begin
                          busy_bit_2 <= _GEN_274;
                        end else if (_T_17) begin
                          busy_bit_2 <= _GEN_210;
                        end else if (_T_39) begin
                          busy_bit_2 <= _GEN_210;
                        end else if (_T_41) begin
                          busy_bit_2 <= _GEN_226;
                        end else begin
                          busy_bit_2 <= _GEN_202;
                        end
                      end else if (_T_49) begin
                        if (3'h2 == io_release_0_rd_addr) begin
                          busy_bit_2 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h2 == io_release_0_rd_addr) begin
                            busy_bit_2 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_2 <= _GEN_210;
                          end else if (_T_39) begin
                            busy_bit_2 <= _GEN_210;
                          end else if (_T_41) begin
                            busy_bit_2 <= _GEN_226;
                          end else begin
                            busy_bit_2 <= _GEN_202;
                          end
                        end else if (_T_44) begin
                          if (3'h2 == io_release_0_rd_addr) begin
                            busy_bit_2 <= 1'h0;
                          end else begin
                            busy_bit_2 <= _GEN_250;
                          end
                        end else if (_T_46) begin
                          busy_bit_2 <= _GEN_274;
                        end else begin
                          busy_bit_2 <= _GEN_250;
                        end
                      end else if (_T_51) begin
                        busy_bit_2 <= _GEN_322;
                      end else if (_T_17) begin
                        busy_bit_2 <= _GEN_258;
                      end else if (_T_44) begin
                        busy_bit_2 <= _GEN_258;
                      end else if (_T_46) begin
                        busy_bit_2 <= _GEN_274;
                      end else begin
                        busy_bit_2 <= _GEN_250;
                      end
                    end else if (_T_54) begin
                      if (3'h2 == io_release_0_rd_addr) begin
                        busy_bit_2 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h2 == io_release_0_rd_addr) begin
                          busy_bit_2 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_2 <= _GEN_258;
                        end else if (_T_44) begin
                          busy_bit_2 <= _GEN_258;
                        end else if (_T_46) begin
                          busy_bit_2 <= _GEN_274;
                        end else begin
                          busy_bit_2 <= _GEN_250;
                        end
                      end else if (_T_49) begin
                        if (3'h2 == io_release_0_rd_addr) begin
                          busy_bit_2 <= 1'h0;
                        end else begin
                          busy_bit_2 <= _GEN_298;
                        end
                      end else if (_T_51) begin
                        busy_bit_2 <= _GEN_322;
                      end else begin
                        busy_bit_2 <= _GEN_298;
                      end
                    end else if (_T_56) begin
                      busy_bit_2 <= _GEN_370;
                    end else if (_T_17) begin
                      busy_bit_2 <= _GEN_306;
                    end else if (_T_49) begin
                      busy_bit_2 <= _GEN_306;
                    end else if (_T_51) begin
                      busy_bit_2 <= _GEN_322;
                    end else begin
                      busy_bit_2 <= _GEN_298;
                    end
                  end else if (_T_21) begin
                    busy_bit_2 <= _GEN_418;
                  end else if (_T_17) begin
                    if (3'h2 == io_release_0_rd_addr) begin
                      busy_bit_2 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_2 <= _GEN_306;
                    end else if (_T_49) begin
                      busy_bit_2 <= _GEN_306;
                    end else if (_T_51) begin
                      busy_bit_2 <= _GEN_322;
                    end else begin
                      busy_bit_2 <= _GEN_298;
                    end
                  end else if (_T_54) begin
                    if (3'h2 == io_release_0_rd_addr) begin
                      busy_bit_2 <= 1'h0;
                    end else begin
                      busy_bit_2 <= _GEN_346;
                    end
                  end else if (_T_56) begin
                    busy_bit_2 <= _GEN_370;
                  end else begin
                    busy_bit_2 <= _GEN_346;
                  end
                end else if (_T_26) begin
                  busy_bit_2 <= _GEN_466;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_2 <= _GEN_354;
                  end else if (_T_54) begin
                    busy_bit_2 <= _GEN_354;
                  end else if (_T_56) begin
                    busy_bit_2 <= _GEN_370;
                  end else begin
                    busy_bit_2 <= _GEN_346;
                  end
                end else if (_T_21) begin
                  busy_bit_2 <= _GEN_418;
                end else if (_T_17) begin
                  busy_bit_2 <= _GEN_354;
                end else if (_T_54) begin
                  busy_bit_2 <= _GEN_354;
                end else if (_T_56) begin
                  busy_bit_2 <= _GEN_370;
                end else begin
                  busy_bit_2 <= _GEN_346;
                end
              end else if (_T_31) begin
                busy_bit_2 <= _GEN_514;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_2 <= _GEN_394;
                end else if (_T_21) begin
                  busy_bit_2 <= _GEN_418;
                end else begin
                  busy_bit_2 <= _GEN_394;
                end
              end else if (_T_26) begin
                busy_bit_2 <= _GEN_466;
              end else if (_T_17) begin
                busy_bit_2 <= _GEN_394;
              end else if (_T_21) begin
                busy_bit_2 <= _GEN_418;
              end else begin
                busy_bit_2 <= _GEN_394;
              end
            end else if (_T_36) begin
              busy_bit_2 <= _GEN_562;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_2 <= _GEN_442;
              end else if (_T_26) begin
                busy_bit_2 <= _GEN_466;
              end else begin
                busy_bit_2 <= _GEN_442;
              end
            end else if (_T_31) begin
              busy_bit_2 <= _GEN_514;
            end else if (_T_17) begin
              busy_bit_2 <= _GEN_442;
            end else if (_T_26) begin
              busy_bit_2 <= _GEN_466;
            end else begin
              busy_bit_2 <= _GEN_442;
            end
          end else if (_T_41) begin
            busy_bit_2 <= _GEN_610;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_2 <= _GEN_490;
            end else if (_T_31) begin
              busy_bit_2 <= _GEN_514;
            end else begin
              busy_bit_2 <= _GEN_490;
            end
          end else if (_T_36) begin
            busy_bit_2 <= _GEN_562;
          end else if (_T_17) begin
            busy_bit_2 <= _GEN_490;
          end else if (_T_31) begin
            busy_bit_2 <= _GEN_514;
          end else begin
            busy_bit_2 <= _GEN_490;
          end
        end else if (_T_46) begin
          busy_bit_2 <= _GEN_658;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_2 <= _GEN_538;
          end else if (_T_36) begin
            busy_bit_2 <= _GEN_562;
          end else begin
            busy_bit_2 <= _GEN_538;
          end
        end else if (_T_41) begin
          busy_bit_2 <= _GEN_610;
        end else if (_T_17) begin
          busy_bit_2 <= _GEN_538;
        end else if (_T_36) begin
          busy_bit_2 <= _GEN_562;
        end else begin
          busy_bit_2 <= _GEN_538;
        end
      end else if (_T_51) begin
        busy_bit_2 <= _GEN_706;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_2 <= _GEN_586;
        end else if (_T_41) begin
          busy_bit_2 <= _GEN_610;
        end else begin
          busy_bit_2 <= _GEN_586;
        end
      end else if (_T_46) begin
        busy_bit_2 <= _GEN_658;
      end else if (_T_17) begin
        busy_bit_2 <= _GEN_586;
      end else if (_T_41) begin
        busy_bit_2 <= _GEN_610;
      end else begin
        busy_bit_2 <= _GEN_586;
      end
    end else if (_T_56) begin
      busy_bit_2 <= _GEN_754;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_2 <= _GEN_634;
      end else if (_T_46) begin
        busy_bit_2 <= _GEN_658;
      end else begin
        busy_bit_2 <= _GEN_634;
      end
    end else if (_T_51) begin
      busy_bit_2 <= _GEN_706;
    end else if (_T_17) begin
      busy_bit_2 <= _GEN_634;
    end else if (_T_46) begin
      busy_bit_2 <= _GEN_658;
    end else begin
      busy_bit_2 <= _GEN_634;
    end
    if (reset) begin
      busy_bit_3 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h3 == io_release_0_rd_addr) begin
                        busy_bit_3 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h3 == io_release_0_rd_addr) begin
                          busy_bit_3 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h3 == io_release_0_rd_addr) begin
                            busy_bit_3 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h3 == io_release_0_rd_addr) begin
                              busy_bit_3 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h3 == io_release_0_rd_addr) begin
                                busy_bit_3 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h3 == io_release_0_rd_addr) begin
                                  busy_bit_3 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h3 == io_release_0_rd_addr) begin
                                    busy_bit_3 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h3 == io_release_0_rd_addr) begin
                                      busy_bit_3 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h3 == io_release_0_rd_addr) begin
                                      busy_bit_3 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_3 <= _GEN_35;
                                  end
                                end else if (_T_24) begin
                                  if (3'h3 == io_release_0_rd_addr) begin
                                    busy_bit_3 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h3 == io_release_0_rd_addr) begin
                                      busy_bit_3 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h3 == io_release_0_rd_addr) begin
                                      busy_bit_3 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_3 <= _GEN_35;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_3 <= _GEN_83;
                                end else if (_T_17) begin
                                  busy_bit_3 <= _GEN_19;
                                end else if (_T_19) begin
                                  busy_bit_3 <= _GEN_19;
                                end else if (_T_21) begin
                                  busy_bit_3 <= _GEN_35;
                                end
                              end else if (_T_29) begin
                                if (3'h3 == io_release_0_rd_addr) begin
                                  busy_bit_3 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h3 == io_release_0_rd_addr) begin
                                    busy_bit_3 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_3 <= _GEN_19;
                                  end else if (_T_19) begin
                                    busy_bit_3 <= _GEN_19;
                                  end else if (_T_21) begin
                                    busy_bit_3 <= _GEN_35;
                                  end
                                end else if (_T_24) begin
                                  if (3'h3 == io_release_0_rd_addr) begin
                                    busy_bit_3 <= 1'h0;
                                  end else begin
                                    busy_bit_3 <= _GEN_59;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_3 <= _GEN_83;
                                end else begin
                                  busy_bit_3 <= _GEN_59;
                                end
                              end else if (_T_31) begin
                                busy_bit_3 <= _GEN_131;
                              end else if (_T_17) begin
                                busy_bit_3 <= _GEN_67;
                              end else if (_T_24) begin
                                busy_bit_3 <= _GEN_67;
                              end else if (_T_26) begin
                                busy_bit_3 <= _GEN_83;
                              end else begin
                                busy_bit_3 <= _GEN_59;
                              end
                            end else if (_T_34) begin
                              if (3'h3 == io_release_0_rd_addr) begin
                                busy_bit_3 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h3 == io_release_0_rd_addr) begin
                                  busy_bit_3 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_3 <= _GEN_67;
                                end else if (_T_24) begin
                                  busy_bit_3 <= _GEN_67;
                                end else if (_T_26) begin
                                  busy_bit_3 <= _GEN_83;
                                end else begin
                                  busy_bit_3 <= _GEN_59;
                                end
                              end else if (_T_29) begin
                                if (3'h3 == io_release_0_rd_addr) begin
                                  busy_bit_3 <= 1'h0;
                                end else begin
                                  busy_bit_3 <= _GEN_107;
                                end
                              end else if (_T_31) begin
                                busy_bit_3 <= _GEN_131;
                              end else begin
                                busy_bit_3 <= _GEN_107;
                              end
                            end else if (_T_36) begin
                              busy_bit_3 <= _GEN_179;
                            end else if (_T_17) begin
                              busy_bit_3 <= _GEN_115;
                            end else if (_T_29) begin
                              busy_bit_3 <= _GEN_115;
                            end else if (_T_31) begin
                              busy_bit_3 <= _GEN_131;
                            end else begin
                              busy_bit_3 <= _GEN_107;
                            end
                          end else if (_T_39) begin
                            if (3'h3 == io_release_0_rd_addr) begin
                              busy_bit_3 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h3 == io_release_0_rd_addr) begin
                                busy_bit_3 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_3 <= _GEN_115;
                              end else if (_T_29) begin
                                busy_bit_3 <= _GEN_115;
                              end else if (_T_31) begin
                                busy_bit_3 <= _GEN_131;
                              end else begin
                                busy_bit_3 <= _GEN_107;
                              end
                            end else if (_T_34) begin
                              if (3'h3 == io_release_0_rd_addr) begin
                                busy_bit_3 <= 1'h0;
                              end else begin
                                busy_bit_3 <= _GEN_155;
                              end
                            end else if (_T_36) begin
                              busy_bit_3 <= _GEN_179;
                            end else begin
                              busy_bit_3 <= _GEN_155;
                            end
                          end else if (_T_41) begin
                            busy_bit_3 <= _GEN_227;
                          end else if (_T_17) begin
                            busy_bit_3 <= _GEN_163;
                          end else if (_T_34) begin
                            busy_bit_3 <= _GEN_163;
                          end else if (_T_36) begin
                            busy_bit_3 <= _GEN_179;
                          end else begin
                            busy_bit_3 <= _GEN_155;
                          end
                        end else if (_T_44) begin
                          if (3'h3 == io_release_0_rd_addr) begin
                            busy_bit_3 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h3 == io_release_0_rd_addr) begin
                              busy_bit_3 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_3 <= _GEN_163;
                            end else if (_T_34) begin
                              busy_bit_3 <= _GEN_163;
                            end else if (_T_36) begin
                              busy_bit_3 <= _GEN_179;
                            end else begin
                              busy_bit_3 <= _GEN_155;
                            end
                          end else if (_T_39) begin
                            if (3'h3 == io_release_0_rd_addr) begin
                              busy_bit_3 <= 1'h0;
                            end else begin
                              busy_bit_3 <= _GEN_203;
                            end
                          end else if (_T_41) begin
                            busy_bit_3 <= _GEN_227;
                          end else begin
                            busy_bit_3 <= _GEN_203;
                          end
                        end else if (_T_46) begin
                          busy_bit_3 <= _GEN_275;
                        end else if (_T_17) begin
                          busy_bit_3 <= _GEN_211;
                        end else if (_T_39) begin
                          busy_bit_3 <= _GEN_211;
                        end else if (_T_41) begin
                          busy_bit_3 <= _GEN_227;
                        end else begin
                          busy_bit_3 <= _GEN_203;
                        end
                      end else if (_T_49) begin
                        if (3'h3 == io_release_0_rd_addr) begin
                          busy_bit_3 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h3 == io_release_0_rd_addr) begin
                            busy_bit_3 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_3 <= _GEN_211;
                          end else if (_T_39) begin
                            busy_bit_3 <= _GEN_211;
                          end else if (_T_41) begin
                            busy_bit_3 <= _GEN_227;
                          end else begin
                            busy_bit_3 <= _GEN_203;
                          end
                        end else if (_T_44) begin
                          if (3'h3 == io_release_0_rd_addr) begin
                            busy_bit_3 <= 1'h0;
                          end else begin
                            busy_bit_3 <= _GEN_251;
                          end
                        end else if (_T_46) begin
                          busy_bit_3 <= _GEN_275;
                        end else begin
                          busy_bit_3 <= _GEN_251;
                        end
                      end else if (_T_51) begin
                        busy_bit_3 <= _GEN_323;
                      end else if (_T_17) begin
                        busy_bit_3 <= _GEN_259;
                      end else if (_T_44) begin
                        busy_bit_3 <= _GEN_259;
                      end else if (_T_46) begin
                        busy_bit_3 <= _GEN_275;
                      end else begin
                        busy_bit_3 <= _GEN_251;
                      end
                    end else if (_T_54) begin
                      if (3'h3 == io_release_0_rd_addr) begin
                        busy_bit_3 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h3 == io_release_0_rd_addr) begin
                          busy_bit_3 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_3 <= _GEN_259;
                        end else if (_T_44) begin
                          busy_bit_3 <= _GEN_259;
                        end else if (_T_46) begin
                          busy_bit_3 <= _GEN_275;
                        end else begin
                          busy_bit_3 <= _GEN_251;
                        end
                      end else if (_T_49) begin
                        if (3'h3 == io_release_0_rd_addr) begin
                          busy_bit_3 <= 1'h0;
                        end else begin
                          busy_bit_3 <= _GEN_299;
                        end
                      end else if (_T_51) begin
                        busy_bit_3 <= _GEN_323;
                      end else begin
                        busy_bit_3 <= _GEN_299;
                      end
                    end else if (_T_56) begin
                      busy_bit_3 <= _GEN_371;
                    end else if (_T_17) begin
                      busy_bit_3 <= _GEN_307;
                    end else if (_T_49) begin
                      busy_bit_3 <= _GEN_307;
                    end else if (_T_51) begin
                      busy_bit_3 <= _GEN_323;
                    end else begin
                      busy_bit_3 <= _GEN_299;
                    end
                  end else if (_T_21) begin
                    busy_bit_3 <= _GEN_419;
                  end else if (_T_17) begin
                    if (3'h3 == io_release_0_rd_addr) begin
                      busy_bit_3 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_3 <= _GEN_307;
                    end else if (_T_49) begin
                      busy_bit_3 <= _GEN_307;
                    end else if (_T_51) begin
                      busy_bit_3 <= _GEN_323;
                    end else begin
                      busy_bit_3 <= _GEN_299;
                    end
                  end else if (_T_54) begin
                    if (3'h3 == io_release_0_rd_addr) begin
                      busy_bit_3 <= 1'h0;
                    end else begin
                      busy_bit_3 <= _GEN_347;
                    end
                  end else if (_T_56) begin
                    busy_bit_3 <= _GEN_371;
                  end else begin
                    busy_bit_3 <= _GEN_347;
                  end
                end else if (_T_26) begin
                  busy_bit_3 <= _GEN_467;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_3 <= _GEN_355;
                  end else if (_T_54) begin
                    busy_bit_3 <= _GEN_355;
                  end else if (_T_56) begin
                    busy_bit_3 <= _GEN_371;
                  end else begin
                    busy_bit_3 <= _GEN_347;
                  end
                end else if (_T_21) begin
                  busy_bit_3 <= _GEN_419;
                end else if (_T_17) begin
                  busy_bit_3 <= _GEN_355;
                end else if (_T_54) begin
                  busy_bit_3 <= _GEN_355;
                end else if (_T_56) begin
                  busy_bit_3 <= _GEN_371;
                end else begin
                  busy_bit_3 <= _GEN_347;
                end
              end else if (_T_31) begin
                busy_bit_3 <= _GEN_515;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_3 <= _GEN_395;
                end else if (_T_21) begin
                  busy_bit_3 <= _GEN_419;
                end else begin
                  busy_bit_3 <= _GEN_395;
                end
              end else if (_T_26) begin
                busy_bit_3 <= _GEN_467;
              end else if (_T_17) begin
                busy_bit_3 <= _GEN_395;
              end else if (_T_21) begin
                busy_bit_3 <= _GEN_419;
              end else begin
                busy_bit_3 <= _GEN_395;
              end
            end else if (_T_36) begin
              busy_bit_3 <= _GEN_563;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_3 <= _GEN_443;
              end else if (_T_26) begin
                busy_bit_3 <= _GEN_467;
              end else begin
                busy_bit_3 <= _GEN_443;
              end
            end else if (_T_31) begin
              busy_bit_3 <= _GEN_515;
            end else if (_T_17) begin
              busy_bit_3 <= _GEN_443;
            end else if (_T_26) begin
              busy_bit_3 <= _GEN_467;
            end else begin
              busy_bit_3 <= _GEN_443;
            end
          end else if (_T_41) begin
            busy_bit_3 <= _GEN_611;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_3 <= _GEN_491;
            end else if (_T_31) begin
              busy_bit_3 <= _GEN_515;
            end else begin
              busy_bit_3 <= _GEN_491;
            end
          end else if (_T_36) begin
            busy_bit_3 <= _GEN_563;
          end else if (_T_17) begin
            busy_bit_3 <= _GEN_491;
          end else if (_T_31) begin
            busy_bit_3 <= _GEN_515;
          end else begin
            busy_bit_3 <= _GEN_491;
          end
        end else if (_T_46) begin
          busy_bit_3 <= _GEN_659;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_3 <= _GEN_539;
          end else if (_T_36) begin
            busy_bit_3 <= _GEN_563;
          end else begin
            busy_bit_3 <= _GEN_539;
          end
        end else if (_T_41) begin
          busy_bit_3 <= _GEN_611;
        end else if (_T_17) begin
          busy_bit_3 <= _GEN_539;
        end else if (_T_36) begin
          busy_bit_3 <= _GEN_563;
        end else begin
          busy_bit_3 <= _GEN_539;
        end
      end else if (_T_51) begin
        busy_bit_3 <= _GEN_707;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_3 <= _GEN_587;
        end else if (_T_41) begin
          busy_bit_3 <= _GEN_611;
        end else begin
          busy_bit_3 <= _GEN_587;
        end
      end else if (_T_46) begin
        busy_bit_3 <= _GEN_659;
      end else if (_T_17) begin
        busy_bit_3 <= _GEN_587;
      end else if (_T_41) begin
        busy_bit_3 <= _GEN_611;
      end else begin
        busy_bit_3 <= _GEN_587;
      end
    end else if (_T_56) begin
      busy_bit_3 <= _GEN_755;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_3 <= _GEN_635;
      end else if (_T_46) begin
        busy_bit_3 <= _GEN_659;
      end else begin
        busy_bit_3 <= _GEN_635;
      end
    end else if (_T_51) begin
      busy_bit_3 <= _GEN_707;
    end else if (_T_17) begin
      busy_bit_3 <= _GEN_635;
    end else if (_T_46) begin
      busy_bit_3 <= _GEN_659;
    end else begin
      busy_bit_3 <= _GEN_635;
    end
    if (reset) begin
      busy_bit_4 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h4 == io_release_0_rd_addr) begin
                        busy_bit_4 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h4 == io_release_0_rd_addr) begin
                          busy_bit_4 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h4 == io_release_0_rd_addr) begin
                            busy_bit_4 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h4 == io_release_0_rd_addr) begin
                              busy_bit_4 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h4 == io_release_0_rd_addr) begin
                                busy_bit_4 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h4 == io_release_0_rd_addr) begin
                                  busy_bit_4 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h4 == io_release_0_rd_addr) begin
                                    busy_bit_4 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h4 == io_release_0_rd_addr) begin
                                      busy_bit_4 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h4 == io_release_0_rd_addr) begin
                                      busy_bit_4 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_4 <= _GEN_36;
                                  end
                                end else if (_T_24) begin
                                  if (3'h4 == io_release_0_rd_addr) begin
                                    busy_bit_4 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h4 == io_release_0_rd_addr) begin
                                      busy_bit_4 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h4 == io_release_0_rd_addr) begin
                                      busy_bit_4 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_4 <= _GEN_36;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_4 <= _GEN_84;
                                end else if (_T_17) begin
                                  busy_bit_4 <= _GEN_20;
                                end else if (_T_19) begin
                                  busy_bit_4 <= _GEN_20;
                                end else if (_T_21) begin
                                  busy_bit_4 <= _GEN_36;
                                end
                              end else if (_T_29) begin
                                if (3'h4 == io_release_0_rd_addr) begin
                                  busy_bit_4 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h4 == io_release_0_rd_addr) begin
                                    busy_bit_4 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_4 <= _GEN_20;
                                  end else if (_T_19) begin
                                    busy_bit_4 <= _GEN_20;
                                  end else if (_T_21) begin
                                    busy_bit_4 <= _GEN_36;
                                  end
                                end else if (_T_24) begin
                                  if (3'h4 == io_release_0_rd_addr) begin
                                    busy_bit_4 <= 1'h0;
                                  end else begin
                                    busy_bit_4 <= _GEN_60;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_4 <= _GEN_84;
                                end else begin
                                  busy_bit_4 <= _GEN_60;
                                end
                              end else if (_T_31) begin
                                busy_bit_4 <= _GEN_132;
                              end else if (_T_17) begin
                                busy_bit_4 <= _GEN_68;
                              end else if (_T_24) begin
                                busy_bit_4 <= _GEN_68;
                              end else if (_T_26) begin
                                busy_bit_4 <= _GEN_84;
                              end else begin
                                busy_bit_4 <= _GEN_60;
                              end
                            end else if (_T_34) begin
                              if (3'h4 == io_release_0_rd_addr) begin
                                busy_bit_4 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h4 == io_release_0_rd_addr) begin
                                  busy_bit_4 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_4 <= _GEN_68;
                                end else if (_T_24) begin
                                  busy_bit_4 <= _GEN_68;
                                end else if (_T_26) begin
                                  busy_bit_4 <= _GEN_84;
                                end else begin
                                  busy_bit_4 <= _GEN_60;
                                end
                              end else if (_T_29) begin
                                if (3'h4 == io_release_0_rd_addr) begin
                                  busy_bit_4 <= 1'h0;
                                end else begin
                                  busy_bit_4 <= _GEN_108;
                                end
                              end else if (_T_31) begin
                                busy_bit_4 <= _GEN_132;
                              end else begin
                                busy_bit_4 <= _GEN_108;
                              end
                            end else if (_T_36) begin
                              busy_bit_4 <= _GEN_180;
                            end else if (_T_17) begin
                              busy_bit_4 <= _GEN_116;
                            end else if (_T_29) begin
                              busy_bit_4 <= _GEN_116;
                            end else if (_T_31) begin
                              busy_bit_4 <= _GEN_132;
                            end else begin
                              busy_bit_4 <= _GEN_108;
                            end
                          end else if (_T_39) begin
                            if (3'h4 == io_release_0_rd_addr) begin
                              busy_bit_4 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h4 == io_release_0_rd_addr) begin
                                busy_bit_4 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_4 <= _GEN_116;
                              end else if (_T_29) begin
                                busy_bit_4 <= _GEN_116;
                              end else if (_T_31) begin
                                busy_bit_4 <= _GEN_132;
                              end else begin
                                busy_bit_4 <= _GEN_108;
                              end
                            end else if (_T_34) begin
                              if (3'h4 == io_release_0_rd_addr) begin
                                busy_bit_4 <= 1'h0;
                              end else begin
                                busy_bit_4 <= _GEN_156;
                              end
                            end else if (_T_36) begin
                              busy_bit_4 <= _GEN_180;
                            end else begin
                              busy_bit_4 <= _GEN_156;
                            end
                          end else if (_T_41) begin
                            busy_bit_4 <= _GEN_228;
                          end else if (_T_17) begin
                            busy_bit_4 <= _GEN_164;
                          end else if (_T_34) begin
                            busy_bit_4 <= _GEN_164;
                          end else if (_T_36) begin
                            busy_bit_4 <= _GEN_180;
                          end else begin
                            busy_bit_4 <= _GEN_156;
                          end
                        end else if (_T_44) begin
                          if (3'h4 == io_release_0_rd_addr) begin
                            busy_bit_4 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h4 == io_release_0_rd_addr) begin
                              busy_bit_4 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_4 <= _GEN_164;
                            end else if (_T_34) begin
                              busy_bit_4 <= _GEN_164;
                            end else if (_T_36) begin
                              busy_bit_4 <= _GEN_180;
                            end else begin
                              busy_bit_4 <= _GEN_156;
                            end
                          end else if (_T_39) begin
                            if (3'h4 == io_release_0_rd_addr) begin
                              busy_bit_4 <= 1'h0;
                            end else begin
                              busy_bit_4 <= _GEN_204;
                            end
                          end else if (_T_41) begin
                            busy_bit_4 <= _GEN_228;
                          end else begin
                            busy_bit_4 <= _GEN_204;
                          end
                        end else if (_T_46) begin
                          busy_bit_4 <= _GEN_276;
                        end else if (_T_17) begin
                          busy_bit_4 <= _GEN_212;
                        end else if (_T_39) begin
                          busy_bit_4 <= _GEN_212;
                        end else if (_T_41) begin
                          busy_bit_4 <= _GEN_228;
                        end else begin
                          busy_bit_4 <= _GEN_204;
                        end
                      end else if (_T_49) begin
                        if (3'h4 == io_release_0_rd_addr) begin
                          busy_bit_4 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h4 == io_release_0_rd_addr) begin
                            busy_bit_4 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_4 <= _GEN_212;
                          end else if (_T_39) begin
                            busy_bit_4 <= _GEN_212;
                          end else if (_T_41) begin
                            busy_bit_4 <= _GEN_228;
                          end else begin
                            busy_bit_4 <= _GEN_204;
                          end
                        end else if (_T_44) begin
                          if (3'h4 == io_release_0_rd_addr) begin
                            busy_bit_4 <= 1'h0;
                          end else begin
                            busy_bit_4 <= _GEN_252;
                          end
                        end else if (_T_46) begin
                          busy_bit_4 <= _GEN_276;
                        end else begin
                          busy_bit_4 <= _GEN_252;
                        end
                      end else if (_T_51) begin
                        busy_bit_4 <= _GEN_324;
                      end else if (_T_17) begin
                        busy_bit_4 <= _GEN_260;
                      end else if (_T_44) begin
                        busy_bit_4 <= _GEN_260;
                      end else if (_T_46) begin
                        busy_bit_4 <= _GEN_276;
                      end else begin
                        busy_bit_4 <= _GEN_252;
                      end
                    end else if (_T_54) begin
                      if (3'h4 == io_release_0_rd_addr) begin
                        busy_bit_4 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h4 == io_release_0_rd_addr) begin
                          busy_bit_4 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_4 <= _GEN_260;
                        end else if (_T_44) begin
                          busy_bit_4 <= _GEN_260;
                        end else if (_T_46) begin
                          busy_bit_4 <= _GEN_276;
                        end else begin
                          busy_bit_4 <= _GEN_252;
                        end
                      end else if (_T_49) begin
                        if (3'h4 == io_release_0_rd_addr) begin
                          busy_bit_4 <= 1'h0;
                        end else begin
                          busy_bit_4 <= _GEN_300;
                        end
                      end else if (_T_51) begin
                        busy_bit_4 <= _GEN_324;
                      end else begin
                        busy_bit_4 <= _GEN_300;
                      end
                    end else if (_T_56) begin
                      busy_bit_4 <= _GEN_372;
                    end else if (_T_17) begin
                      busy_bit_4 <= _GEN_308;
                    end else if (_T_49) begin
                      busy_bit_4 <= _GEN_308;
                    end else if (_T_51) begin
                      busy_bit_4 <= _GEN_324;
                    end else begin
                      busy_bit_4 <= _GEN_300;
                    end
                  end else if (_T_21) begin
                    busy_bit_4 <= _GEN_420;
                  end else if (_T_17) begin
                    if (3'h4 == io_release_0_rd_addr) begin
                      busy_bit_4 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_4 <= _GEN_308;
                    end else if (_T_49) begin
                      busy_bit_4 <= _GEN_308;
                    end else if (_T_51) begin
                      busy_bit_4 <= _GEN_324;
                    end else begin
                      busy_bit_4 <= _GEN_300;
                    end
                  end else if (_T_54) begin
                    if (3'h4 == io_release_0_rd_addr) begin
                      busy_bit_4 <= 1'h0;
                    end else begin
                      busy_bit_4 <= _GEN_348;
                    end
                  end else if (_T_56) begin
                    busy_bit_4 <= _GEN_372;
                  end else begin
                    busy_bit_4 <= _GEN_348;
                  end
                end else if (_T_26) begin
                  busy_bit_4 <= _GEN_468;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_4 <= _GEN_356;
                  end else if (_T_54) begin
                    busy_bit_4 <= _GEN_356;
                  end else if (_T_56) begin
                    busy_bit_4 <= _GEN_372;
                  end else begin
                    busy_bit_4 <= _GEN_348;
                  end
                end else if (_T_21) begin
                  busy_bit_4 <= _GEN_420;
                end else if (_T_17) begin
                  busy_bit_4 <= _GEN_356;
                end else if (_T_54) begin
                  busy_bit_4 <= _GEN_356;
                end else if (_T_56) begin
                  busy_bit_4 <= _GEN_372;
                end else begin
                  busy_bit_4 <= _GEN_348;
                end
              end else if (_T_31) begin
                busy_bit_4 <= _GEN_516;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_4 <= _GEN_396;
                end else if (_T_21) begin
                  busy_bit_4 <= _GEN_420;
                end else begin
                  busy_bit_4 <= _GEN_396;
                end
              end else if (_T_26) begin
                busy_bit_4 <= _GEN_468;
              end else if (_T_17) begin
                busy_bit_4 <= _GEN_396;
              end else if (_T_21) begin
                busy_bit_4 <= _GEN_420;
              end else begin
                busy_bit_4 <= _GEN_396;
              end
            end else if (_T_36) begin
              busy_bit_4 <= _GEN_564;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_4 <= _GEN_444;
              end else if (_T_26) begin
                busy_bit_4 <= _GEN_468;
              end else begin
                busy_bit_4 <= _GEN_444;
              end
            end else if (_T_31) begin
              busy_bit_4 <= _GEN_516;
            end else if (_T_17) begin
              busy_bit_4 <= _GEN_444;
            end else if (_T_26) begin
              busy_bit_4 <= _GEN_468;
            end else begin
              busy_bit_4 <= _GEN_444;
            end
          end else if (_T_41) begin
            busy_bit_4 <= _GEN_612;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_4 <= _GEN_492;
            end else if (_T_31) begin
              busy_bit_4 <= _GEN_516;
            end else begin
              busy_bit_4 <= _GEN_492;
            end
          end else if (_T_36) begin
            busy_bit_4 <= _GEN_564;
          end else if (_T_17) begin
            busy_bit_4 <= _GEN_492;
          end else if (_T_31) begin
            busy_bit_4 <= _GEN_516;
          end else begin
            busy_bit_4 <= _GEN_492;
          end
        end else if (_T_46) begin
          busy_bit_4 <= _GEN_660;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_4 <= _GEN_540;
          end else if (_T_36) begin
            busy_bit_4 <= _GEN_564;
          end else begin
            busy_bit_4 <= _GEN_540;
          end
        end else if (_T_41) begin
          busy_bit_4 <= _GEN_612;
        end else if (_T_17) begin
          busy_bit_4 <= _GEN_540;
        end else if (_T_36) begin
          busy_bit_4 <= _GEN_564;
        end else begin
          busy_bit_4 <= _GEN_540;
        end
      end else if (_T_51) begin
        busy_bit_4 <= _GEN_708;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_4 <= _GEN_588;
        end else if (_T_41) begin
          busy_bit_4 <= _GEN_612;
        end else begin
          busy_bit_4 <= _GEN_588;
        end
      end else if (_T_46) begin
        busy_bit_4 <= _GEN_660;
      end else if (_T_17) begin
        busy_bit_4 <= _GEN_588;
      end else if (_T_41) begin
        busy_bit_4 <= _GEN_612;
      end else begin
        busy_bit_4 <= _GEN_588;
      end
    end else if (_T_56) begin
      busy_bit_4 <= _GEN_756;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_4 <= _GEN_636;
      end else if (_T_46) begin
        busy_bit_4 <= _GEN_660;
      end else begin
        busy_bit_4 <= _GEN_636;
      end
    end else if (_T_51) begin
      busy_bit_4 <= _GEN_708;
    end else if (_T_17) begin
      busy_bit_4 <= _GEN_636;
    end else if (_T_46) begin
      busy_bit_4 <= _GEN_660;
    end else begin
      busy_bit_4 <= _GEN_636;
    end
    if (reset) begin
      busy_bit_5 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h5 == io_release_0_rd_addr) begin
                        busy_bit_5 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h5 == io_release_0_rd_addr) begin
                          busy_bit_5 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h5 == io_release_0_rd_addr) begin
                            busy_bit_5 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h5 == io_release_0_rd_addr) begin
                              busy_bit_5 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h5 == io_release_0_rd_addr) begin
                                busy_bit_5 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h5 == io_release_0_rd_addr) begin
                                  busy_bit_5 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h5 == io_release_0_rd_addr) begin
                                    busy_bit_5 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h5 == io_release_0_rd_addr) begin
                                      busy_bit_5 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h5 == io_release_0_rd_addr) begin
                                      busy_bit_5 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_5 <= _GEN_37;
                                  end
                                end else if (_T_24) begin
                                  if (3'h5 == io_release_0_rd_addr) begin
                                    busy_bit_5 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h5 == io_release_0_rd_addr) begin
                                      busy_bit_5 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h5 == io_release_0_rd_addr) begin
                                      busy_bit_5 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_5 <= _GEN_37;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_5 <= _GEN_85;
                                end else if (_T_17) begin
                                  busy_bit_5 <= _GEN_21;
                                end else if (_T_19) begin
                                  busy_bit_5 <= _GEN_21;
                                end else if (_T_21) begin
                                  busy_bit_5 <= _GEN_37;
                                end
                              end else if (_T_29) begin
                                if (3'h5 == io_release_0_rd_addr) begin
                                  busy_bit_5 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h5 == io_release_0_rd_addr) begin
                                    busy_bit_5 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_5 <= _GEN_21;
                                  end else if (_T_19) begin
                                    busy_bit_5 <= _GEN_21;
                                  end else if (_T_21) begin
                                    busy_bit_5 <= _GEN_37;
                                  end
                                end else if (_T_24) begin
                                  if (3'h5 == io_release_0_rd_addr) begin
                                    busy_bit_5 <= 1'h0;
                                  end else begin
                                    busy_bit_5 <= _GEN_61;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_5 <= _GEN_85;
                                end else begin
                                  busy_bit_5 <= _GEN_61;
                                end
                              end else if (_T_31) begin
                                busy_bit_5 <= _GEN_133;
                              end else if (_T_17) begin
                                busy_bit_5 <= _GEN_69;
                              end else if (_T_24) begin
                                busy_bit_5 <= _GEN_69;
                              end else if (_T_26) begin
                                busy_bit_5 <= _GEN_85;
                              end else begin
                                busy_bit_5 <= _GEN_61;
                              end
                            end else if (_T_34) begin
                              if (3'h5 == io_release_0_rd_addr) begin
                                busy_bit_5 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h5 == io_release_0_rd_addr) begin
                                  busy_bit_5 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_5 <= _GEN_69;
                                end else if (_T_24) begin
                                  busy_bit_5 <= _GEN_69;
                                end else if (_T_26) begin
                                  busy_bit_5 <= _GEN_85;
                                end else begin
                                  busy_bit_5 <= _GEN_61;
                                end
                              end else if (_T_29) begin
                                if (3'h5 == io_release_0_rd_addr) begin
                                  busy_bit_5 <= 1'h0;
                                end else begin
                                  busy_bit_5 <= _GEN_109;
                                end
                              end else if (_T_31) begin
                                busy_bit_5 <= _GEN_133;
                              end else begin
                                busy_bit_5 <= _GEN_109;
                              end
                            end else if (_T_36) begin
                              busy_bit_5 <= _GEN_181;
                            end else if (_T_17) begin
                              busy_bit_5 <= _GEN_117;
                            end else if (_T_29) begin
                              busy_bit_5 <= _GEN_117;
                            end else if (_T_31) begin
                              busy_bit_5 <= _GEN_133;
                            end else begin
                              busy_bit_5 <= _GEN_109;
                            end
                          end else if (_T_39) begin
                            if (3'h5 == io_release_0_rd_addr) begin
                              busy_bit_5 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h5 == io_release_0_rd_addr) begin
                                busy_bit_5 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_5 <= _GEN_117;
                              end else if (_T_29) begin
                                busy_bit_5 <= _GEN_117;
                              end else if (_T_31) begin
                                busy_bit_5 <= _GEN_133;
                              end else begin
                                busy_bit_5 <= _GEN_109;
                              end
                            end else if (_T_34) begin
                              if (3'h5 == io_release_0_rd_addr) begin
                                busy_bit_5 <= 1'h0;
                              end else begin
                                busy_bit_5 <= _GEN_157;
                              end
                            end else if (_T_36) begin
                              busy_bit_5 <= _GEN_181;
                            end else begin
                              busy_bit_5 <= _GEN_157;
                            end
                          end else if (_T_41) begin
                            busy_bit_5 <= _GEN_229;
                          end else if (_T_17) begin
                            busy_bit_5 <= _GEN_165;
                          end else if (_T_34) begin
                            busy_bit_5 <= _GEN_165;
                          end else if (_T_36) begin
                            busy_bit_5 <= _GEN_181;
                          end else begin
                            busy_bit_5 <= _GEN_157;
                          end
                        end else if (_T_44) begin
                          if (3'h5 == io_release_0_rd_addr) begin
                            busy_bit_5 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h5 == io_release_0_rd_addr) begin
                              busy_bit_5 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_5 <= _GEN_165;
                            end else if (_T_34) begin
                              busy_bit_5 <= _GEN_165;
                            end else if (_T_36) begin
                              busy_bit_5 <= _GEN_181;
                            end else begin
                              busy_bit_5 <= _GEN_157;
                            end
                          end else if (_T_39) begin
                            if (3'h5 == io_release_0_rd_addr) begin
                              busy_bit_5 <= 1'h0;
                            end else begin
                              busy_bit_5 <= _GEN_205;
                            end
                          end else if (_T_41) begin
                            busy_bit_5 <= _GEN_229;
                          end else begin
                            busy_bit_5 <= _GEN_205;
                          end
                        end else if (_T_46) begin
                          busy_bit_5 <= _GEN_277;
                        end else if (_T_17) begin
                          busy_bit_5 <= _GEN_213;
                        end else if (_T_39) begin
                          busy_bit_5 <= _GEN_213;
                        end else if (_T_41) begin
                          busy_bit_5 <= _GEN_229;
                        end else begin
                          busy_bit_5 <= _GEN_205;
                        end
                      end else if (_T_49) begin
                        if (3'h5 == io_release_0_rd_addr) begin
                          busy_bit_5 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h5 == io_release_0_rd_addr) begin
                            busy_bit_5 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_5 <= _GEN_213;
                          end else if (_T_39) begin
                            busy_bit_5 <= _GEN_213;
                          end else if (_T_41) begin
                            busy_bit_5 <= _GEN_229;
                          end else begin
                            busy_bit_5 <= _GEN_205;
                          end
                        end else if (_T_44) begin
                          if (3'h5 == io_release_0_rd_addr) begin
                            busy_bit_5 <= 1'h0;
                          end else begin
                            busy_bit_5 <= _GEN_253;
                          end
                        end else if (_T_46) begin
                          busy_bit_5 <= _GEN_277;
                        end else begin
                          busy_bit_5 <= _GEN_253;
                        end
                      end else if (_T_51) begin
                        busy_bit_5 <= _GEN_325;
                      end else if (_T_17) begin
                        busy_bit_5 <= _GEN_261;
                      end else if (_T_44) begin
                        busy_bit_5 <= _GEN_261;
                      end else if (_T_46) begin
                        busy_bit_5 <= _GEN_277;
                      end else begin
                        busy_bit_5 <= _GEN_253;
                      end
                    end else if (_T_54) begin
                      if (3'h5 == io_release_0_rd_addr) begin
                        busy_bit_5 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h5 == io_release_0_rd_addr) begin
                          busy_bit_5 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_5 <= _GEN_261;
                        end else if (_T_44) begin
                          busy_bit_5 <= _GEN_261;
                        end else if (_T_46) begin
                          busy_bit_5 <= _GEN_277;
                        end else begin
                          busy_bit_5 <= _GEN_253;
                        end
                      end else if (_T_49) begin
                        if (3'h5 == io_release_0_rd_addr) begin
                          busy_bit_5 <= 1'h0;
                        end else begin
                          busy_bit_5 <= _GEN_301;
                        end
                      end else if (_T_51) begin
                        busy_bit_5 <= _GEN_325;
                      end else begin
                        busy_bit_5 <= _GEN_301;
                      end
                    end else if (_T_56) begin
                      busy_bit_5 <= _GEN_373;
                    end else if (_T_17) begin
                      busy_bit_5 <= _GEN_309;
                    end else if (_T_49) begin
                      busy_bit_5 <= _GEN_309;
                    end else if (_T_51) begin
                      busy_bit_5 <= _GEN_325;
                    end else begin
                      busy_bit_5 <= _GEN_301;
                    end
                  end else if (_T_21) begin
                    busy_bit_5 <= _GEN_421;
                  end else if (_T_17) begin
                    if (3'h5 == io_release_0_rd_addr) begin
                      busy_bit_5 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_5 <= _GEN_309;
                    end else if (_T_49) begin
                      busy_bit_5 <= _GEN_309;
                    end else if (_T_51) begin
                      busy_bit_5 <= _GEN_325;
                    end else begin
                      busy_bit_5 <= _GEN_301;
                    end
                  end else if (_T_54) begin
                    if (3'h5 == io_release_0_rd_addr) begin
                      busy_bit_5 <= 1'h0;
                    end else begin
                      busy_bit_5 <= _GEN_349;
                    end
                  end else if (_T_56) begin
                    busy_bit_5 <= _GEN_373;
                  end else begin
                    busy_bit_5 <= _GEN_349;
                  end
                end else if (_T_26) begin
                  busy_bit_5 <= _GEN_469;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_5 <= _GEN_357;
                  end else if (_T_54) begin
                    busy_bit_5 <= _GEN_357;
                  end else if (_T_56) begin
                    busy_bit_5 <= _GEN_373;
                  end else begin
                    busy_bit_5 <= _GEN_349;
                  end
                end else if (_T_21) begin
                  busy_bit_5 <= _GEN_421;
                end else if (_T_17) begin
                  busy_bit_5 <= _GEN_357;
                end else if (_T_54) begin
                  busy_bit_5 <= _GEN_357;
                end else if (_T_56) begin
                  busy_bit_5 <= _GEN_373;
                end else begin
                  busy_bit_5 <= _GEN_349;
                end
              end else if (_T_31) begin
                busy_bit_5 <= _GEN_517;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_5 <= _GEN_397;
                end else if (_T_21) begin
                  busy_bit_5 <= _GEN_421;
                end else begin
                  busy_bit_5 <= _GEN_397;
                end
              end else if (_T_26) begin
                busy_bit_5 <= _GEN_469;
              end else if (_T_17) begin
                busy_bit_5 <= _GEN_397;
              end else if (_T_21) begin
                busy_bit_5 <= _GEN_421;
              end else begin
                busy_bit_5 <= _GEN_397;
              end
            end else if (_T_36) begin
              busy_bit_5 <= _GEN_565;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_5 <= _GEN_445;
              end else if (_T_26) begin
                busy_bit_5 <= _GEN_469;
              end else begin
                busy_bit_5 <= _GEN_445;
              end
            end else if (_T_31) begin
              busy_bit_5 <= _GEN_517;
            end else if (_T_17) begin
              busy_bit_5 <= _GEN_445;
            end else if (_T_26) begin
              busy_bit_5 <= _GEN_469;
            end else begin
              busy_bit_5 <= _GEN_445;
            end
          end else if (_T_41) begin
            busy_bit_5 <= _GEN_613;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_5 <= _GEN_493;
            end else if (_T_31) begin
              busy_bit_5 <= _GEN_517;
            end else begin
              busy_bit_5 <= _GEN_493;
            end
          end else if (_T_36) begin
            busy_bit_5 <= _GEN_565;
          end else if (_T_17) begin
            busy_bit_5 <= _GEN_493;
          end else if (_T_31) begin
            busy_bit_5 <= _GEN_517;
          end else begin
            busy_bit_5 <= _GEN_493;
          end
        end else if (_T_46) begin
          busy_bit_5 <= _GEN_661;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_5 <= _GEN_541;
          end else if (_T_36) begin
            busy_bit_5 <= _GEN_565;
          end else begin
            busy_bit_5 <= _GEN_541;
          end
        end else if (_T_41) begin
          busy_bit_5 <= _GEN_613;
        end else if (_T_17) begin
          busy_bit_5 <= _GEN_541;
        end else if (_T_36) begin
          busy_bit_5 <= _GEN_565;
        end else begin
          busy_bit_5 <= _GEN_541;
        end
      end else if (_T_51) begin
        busy_bit_5 <= _GEN_709;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_5 <= _GEN_589;
        end else if (_T_41) begin
          busy_bit_5 <= _GEN_613;
        end else begin
          busy_bit_5 <= _GEN_589;
        end
      end else if (_T_46) begin
        busy_bit_5 <= _GEN_661;
      end else if (_T_17) begin
        busy_bit_5 <= _GEN_589;
      end else if (_T_41) begin
        busy_bit_5 <= _GEN_613;
      end else begin
        busy_bit_5 <= _GEN_589;
      end
    end else if (_T_56) begin
      busy_bit_5 <= _GEN_757;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_5 <= _GEN_637;
      end else if (_T_46) begin
        busy_bit_5 <= _GEN_661;
      end else begin
        busy_bit_5 <= _GEN_637;
      end
    end else if (_T_51) begin
      busy_bit_5 <= _GEN_709;
    end else if (_T_17) begin
      busy_bit_5 <= _GEN_637;
    end else if (_T_46) begin
      busy_bit_5 <= _GEN_661;
    end else begin
      busy_bit_5 <= _GEN_637;
    end
    if (reset) begin
      busy_bit_6 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h6 == io_release_0_rd_addr) begin
                        busy_bit_6 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h6 == io_release_0_rd_addr) begin
                          busy_bit_6 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h6 == io_release_0_rd_addr) begin
                            busy_bit_6 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h6 == io_release_0_rd_addr) begin
                              busy_bit_6 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h6 == io_release_0_rd_addr) begin
                                busy_bit_6 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h6 == io_release_0_rd_addr) begin
                                  busy_bit_6 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h6 == io_release_0_rd_addr) begin
                                    busy_bit_6 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h6 == io_release_0_rd_addr) begin
                                      busy_bit_6 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h6 == io_release_0_rd_addr) begin
                                      busy_bit_6 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_6 <= _GEN_38;
                                  end
                                end else if (_T_24) begin
                                  if (3'h6 == io_release_0_rd_addr) begin
                                    busy_bit_6 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h6 == io_release_0_rd_addr) begin
                                      busy_bit_6 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h6 == io_release_0_rd_addr) begin
                                      busy_bit_6 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_6 <= _GEN_38;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_6 <= _GEN_86;
                                end else if (_T_17) begin
                                  busy_bit_6 <= _GEN_22;
                                end else if (_T_19) begin
                                  busy_bit_6 <= _GEN_22;
                                end else if (_T_21) begin
                                  busy_bit_6 <= _GEN_38;
                                end
                              end else if (_T_29) begin
                                if (3'h6 == io_release_0_rd_addr) begin
                                  busy_bit_6 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h6 == io_release_0_rd_addr) begin
                                    busy_bit_6 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_6 <= _GEN_22;
                                  end else if (_T_19) begin
                                    busy_bit_6 <= _GEN_22;
                                  end else if (_T_21) begin
                                    busy_bit_6 <= _GEN_38;
                                  end
                                end else if (_T_24) begin
                                  if (3'h6 == io_release_0_rd_addr) begin
                                    busy_bit_6 <= 1'h0;
                                  end else begin
                                    busy_bit_6 <= _GEN_62;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_6 <= _GEN_86;
                                end else begin
                                  busy_bit_6 <= _GEN_62;
                                end
                              end else if (_T_31) begin
                                busy_bit_6 <= _GEN_134;
                              end else if (_T_17) begin
                                busy_bit_6 <= _GEN_70;
                              end else if (_T_24) begin
                                busy_bit_6 <= _GEN_70;
                              end else if (_T_26) begin
                                busy_bit_6 <= _GEN_86;
                              end else begin
                                busy_bit_6 <= _GEN_62;
                              end
                            end else if (_T_34) begin
                              if (3'h6 == io_release_0_rd_addr) begin
                                busy_bit_6 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h6 == io_release_0_rd_addr) begin
                                  busy_bit_6 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_6 <= _GEN_70;
                                end else if (_T_24) begin
                                  busy_bit_6 <= _GEN_70;
                                end else if (_T_26) begin
                                  busy_bit_6 <= _GEN_86;
                                end else begin
                                  busy_bit_6 <= _GEN_62;
                                end
                              end else if (_T_29) begin
                                if (3'h6 == io_release_0_rd_addr) begin
                                  busy_bit_6 <= 1'h0;
                                end else begin
                                  busy_bit_6 <= _GEN_110;
                                end
                              end else if (_T_31) begin
                                busy_bit_6 <= _GEN_134;
                              end else begin
                                busy_bit_6 <= _GEN_110;
                              end
                            end else if (_T_36) begin
                              busy_bit_6 <= _GEN_182;
                            end else if (_T_17) begin
                              busy_bit_6 <= _GEN_118;
                            end else if (_T_29) begin
                              busy_bit_6 <= _GEN_118;
                            end else if (_T_31) begin
                              busy_bit_6 <= _GEN_134;
                            end else begin
                              busy_bit_6 <= _GEN_110;
                            end
                          end else if (_T_39) begin
                            if (3'h6 == io_release_0_rd_addr) begin
                              busy_bit_6 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h6 == io_release_0_rd_addr) begin
                                busy_bit_6 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_6 <= _GEN_118;
                              end else if (_T_29) begin
                                busy_bit_6 <= _GEN_118;
                              end else if (_T_31) begin
                                busy_bit_6 <= _GEN_134;
                              end else begin
                                busy_bit_6 <= _GEN_110;
                              end
                            end else if (_T_34) begin
                              if (3'h6 == io_release_0_rd_addr) begin
                                busy_bit_6 <= 1'h0;
                              end else begin
                                busy_bit_6 <= _GEN_158;
                              end
                            end else if (_T_36) begin
                              busy_bit_6 <= _GEN_182;
                            end else begin
                              busy_bit_6 <= _GEN_158;
                            end
                          end else if (_T_41) begin
                            busy_bit_6 <= _GEN_230;
                          end else if (_T_17) begin
                            busy_bit_6 <= _GEN_166;
                          end else if (_T_34) begin
                            busy_bit_6 <= _GEN_166;
                          end else if (_T_36) begin
                            busy_bit_6 <= _GEN_182;
                          end else begin
                            busy_bit_6 <= _GEN_158;
                          end
                        end else if (_T_44) begin
                          if (3'h6 == io_release_0_rd_addr) begin
                            busy_bit_6 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h6 == io_release_0_rd_addr) begin
                              busy_bit_6 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_6 <= _GEN_166;
                            end else if (_T_34) begin
                              busy_bit_6 <= _GEN_166;
                            end else if (_T_36) begin
                              busy_bit_6 <= _GEN_182;
                            end else begin
                              busy_bit_6 <= _GEN_158;
                            end
                          end else if (_T_39) begin
                            if (3'h6 == io_release_0_rd_addr) begin
                              busy_bit_6 <= 1'h0;
                            end else begin
                              busy_bit_6 <= _GEN_206;
                            end
                          end else if (_T_41) begin
                            busy_bit_6 <= _GEN_230;
                          end else begin
                            busy_bit_6 <= _GEN_206;
                          end
                        end else if (_T_46) begin
                          busy_bit_6 <= _GEN_278;
                        end else if (_T_17) begin
                          busy_bit_6 <= _GEN_214;
                        end else if (_T_39) begin
                          busy_bit_6 <= _GEN_214;
                        end else if (_T_41) begin
                          busy_bit_6 <= _GEN_230;
                        end else begin
                          busy_bit_6 <= _GEN_206;
                        end
                      end else if (_T_49) begin
                        if (3'h6 == io_release_0_rd_addr) begin
                          busy_bit_6 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h6 == io_release_0_rd_addr) begin
                            busy_bit_6 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_6 <= _GEN_214;
                          end else if (_T_39) begin
                            busy_bit_6 <= _GEN_214;
                          end else if (_T_41) begin
                            busy_bit_6 <= _GEN_230;
                          end else begin
                            busy_bit_6 <= _GEN_206;
                          end
                        end else if (_T_44) begin
                          if (3'h6 == io_release_0_rd_addr) begin
                            busy_bit_6 <= 1'h0;
                          end else begin
                            busy_bit_6 <= _GEN_254;
                          end
                        end else if (_T_46) begin
                          busy_bit_6 <= _GEN_278;
                        end else begin
                          busy_bit_6 <= _GEN_254;
                        end
                      end else if (_T_51) begin
                        busy_bit_6 <= _GEN_326;
                      end else if (_T_17) begin
                        busy_bit_6 <= _GEN_262;
                      end else if (_T_44) begin
                        busy_bit_6 <= _GEN_262;
                      end else if (_T_46) begin
                        busy_bit_6 <= _GEN_278;
                      end else begin
                        busy_bit_6 <= _GEN_254;
                      end
                    end else if (_T_54) begin
                      if (3'h6 == io_release_0_rd_addr) begin
                        busy_bit_6 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h6 == io_release_0_rd_addr) begin
                          busy_bit_6 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_6 <= _GEN_262;
                        end else if (_T_44) begin
                          busy_bit_6 <= _GEN_262;
                        end else if (_T_46) begin
                          busy_bit_6 <= _GEN_278;
                        end else begin
                          busy_bit_6 <= _GEN_254;
                        end
                      end else if (_T_49) begin
                        if (3'h6 == io_release_0_rd_addr) begin
                          busy_bit_6 <= 1'h0;
                        end else begin
                          busy_bit_6 <= _GEN_302;
                        end
                      end else if (_T_51) begin
                        busy_bit_6 <= _GEN_326;
                      end else begin
                        busy_bit_6 <= _GEN_302;
                      end
                    end else if (_T_56) begin
                      busy_bit_6 <= _GEN_374;
                    end else if (_T_17) begin
                      busy_bit_6 <= _GEN_310;
                    end else if (_T_49) begin
                      busy_bit_6 <= _GEN_310;
                    end else if (_T_51) begin
                      busy_bit_6 <= _GEN_326;
                    end else begin
                      busy_bit_6 <= _GEN_302;
                    end
                  end else if (_T_21) begin
                    busy_bit_6 <= _GEN_422;
                  end else if (_T_17) begin
                    if (3'h6 == io_release_0_rd_addr) begin
                      busy_bit_6 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_6 <= _GEN_310;
                    end else if (_T_49) begin
                      busy_bit_6 <= _GEN_310;
                    end else if (_T_51) begin
                      busy_bit_6 <= _GEN_326;
                    end else begin
                      busy_bit_6 <= _GEN_302;
                    end
                  end else if (_T_54) begin
                    if (3'h6 == io_release_0_rd_addr) begin
                      busy_bit_6 <= 1'h0;
                    end else begin
                      busy_bit_6 <= _GEN_350;
                    end
                  end else if (_T_56) begin
                    busy_bit_6 <= _GEN_374;
                  end else begin
                    busy_bit_6 <= _GEN_350;
                  end
                end else if (_T_26) begin
                  busy_bit_6 <= _GEN_470;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_6 <= _GEN_358;
                  end else if (_T_54) begin
                    busy_bit_6 <= _GEN_358;
                  end else if (_T_56) begin
                    busy_bit_6 <= _GEN_374;
                  end else begin
                    busy_bit_6 <= _GEN_350;
                  end
                end else if (_T_21) begin
                  busy_bit_6 <= _GEN_422;
                end else if (_T_17) begin
                  busy_bit_6 <= _GEN_358;
                end else if (_T_54) begin
                  busy_bit_6 <= _GEN_358;
                end else if (_T_56) begin
                  busy_bit_6 <= _GEN_374;
                end else begin
                  busy_bit_6 <= _GEN_350;
                end
              end else if (_T_31) begin
                busy_bit_6 <= _GEN_518;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_6 <= _GEN_398;
                end else if (_T_21) begin
                  busy_bit_6 <= _GEN_422;
                end else begin
                  busy_bit_6 <= _GEN_398;
                end
              end else if (_T_26) begin
                busy_bit_6 <= _GEN_470;
              end else if (_T_17) begin
                busy_bit_6 <= _GEN_398;
              end else if (_T_21) begin
                busy_bit_6 <= _GEN_422;
              end else begin
                busy_bit_6 <= _GEN_398;
              end
            end else if (_T_36) begin
              busy_bit_6 <= _GEN_566;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_6 <= _GEN_446;
              end else if (_T_26) begin
                busy_bit_6 <= _GEN_470;
              end else begin
                busy_bit_6 <= _GEN_446;
              end
            end else if (_T_31) begin
              busy_bit_6 <= _GEN_518;
            end else if (_T_17) begin
              busy_bit_6 <= _GEN_446;
            end else if (_T_26) begin
              busy_bit_6 <= _GEN_470;
            end else begin
              busy_bit_6 <= _GEN_446;
            end
          end else if (_T_41) begin
            busy_bit_6 <= _GEN_614;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_6 <= _GEN_494;
            end else if (_T_31) begin
              busy_bit_6 <= _GEN_518;
            end else begin
              busy_bit_6 <= _GEN_494;
            end
          end else if (_T_36) begin
            busy_bit_6 <= _GEN_566;
          end else if (_T_17) begin
            busy_bit_6 <= _GEN_494;
          end else if (_T_31) begin
            busy_bit_6 <= _GEN_518;
          end else begin
            busy_bit_6 <= _GEN_494;
          end
        end else if (_T_46) begin
          busy_bit_6 <= _GEN_662;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_6 <= _GEN_542;
          end else if (_T_36) begin
            busy_bit_6 <= _GEN_566;
          end else begin
            busy_bit_6 <= _GEN_542;
          end
        end else if (_T_41) begin
          busy_bit_6 <= _GEN_614;
        end else if (_T_17) begin
          busy_bit_6 <= _GEN_542;
        end else if (_T_36) begin
          busy_bit_6 <= _GEN_566;
        end else begin
          busy_bit_6 <= _GEN_542;
        end
      end else if (_T_51) begin
        busy_bit_6 <= _GEN_710;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_6 <= _GEN_590;
        end else if (_T_41) begin
          busy_bit_6 <= _GEN_614;
        end else begin
          busy_bit_6 <= _GEN_590;
        end
      end else if (_T_46) begin
        busy_bit_6 <= _GEN_662;
      end else if (_T_17) begin
        busy_bit_6 <= _GEN_590;
      end else if (_T_41) begin
        busy_bit_6 <= _GEN_614;
      end else begin
        busy_bit_6 <= _GEN_590;
      end
    end else if (_T_56) begin
      busy_bit_6 <= _GEN_758;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_6 <= _GEN_638;
      end else if (_T_46) begin
        busy_bit_6 <= _GEN_662;
      end else begin
        busy_bit_6 <= _GEN_638;
      end
    end else if (_T_51) begin
      busy_bit_6 <= _GEN_710;
    end else if (_T_17) begin
      busy_bit_6 <= _GEN_638;
    end else if (_T_46) begin
      busy_bit_6 <= _GEN_662;
    end else begin
      busy_bit_6 <= _GEN_638;
    end
    if (reset) begin
      busy_bit_7 <= 1'h0;
    end else if (_T_17) begin
      if (_T_17) begin
        if (_T_17) begin
          if (_T_17) begin
            if (_T_17) begin
              if (_T_17) begin
                if (_T_17) begin
                  if (_T_17) begin
                    if (_T_17) begin
                      if (3'h7 == io_release_0_rd_addr) begin
                        busy_bit_7 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h7 == io_release_0_rd_addr) begin
                          busy_bit_7 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h7 == io_release_0_rd_addr) begin
                            busy_bit_7 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h7 == io_release_0_rd_addr) begin
                              busy_bit_7 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h7 == io_release_0_rd_addr) begin
                                busy_bit_7 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h7 == io_release_0_rd_addr) begin
                                  busy_bit_7 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h7 == io_release_0_rd_addr) begin
                                    busy_bit_7 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h7 == io_release_0_rd_addr) begin
                                      busy_bit_7 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h7 == io_release_0_rd_addr) begin
                                      busy_bit_7 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_7 <= _GEN_39;
                                  end
                                end else if (_T_24) begin
                                  if (3'h7 == io_release_0_rd_addr) begin
                                    busy_bit_7 <= 1'h0;
                                  end else if (_T_17) begin
                                    if (3'h7 == io_release_0_rd_addr) begin
                                      busy_bit_7 <= 1'h0;
                                    end
                                  end else if (_T_19) begin
                                    if (3'h7 == io_release_0_rd_addr) begin
                                      busy_bit_7 <= 1'h0;
                                    end
                                  end else if (_T_21) begin
                                    busy_bit_7 <= _GEN_39;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_7 <= _GEN_87;
                                end else if (_T_17) begin
                                  busy_bit_7 <= _GEN_23;
                                end else if (_T_19) begin
                                  busy_bit_7 <= _GEN_23;
                                end else if (_T_21) begin
                                  busy_bit_7 <= _GEN_39;
                                end
                              end else if (_T_29) begin
                                if (3'h7 == io_release_0_rd_addr) begin
                                  busy_bit_7 <= 1'h0;
                                end else if (_T_17) begin
                                  if (3'h7 == io_release_0_rd_addr) begin
                                    busy_bit_7 <= 1'h0;
                                  end else if (_T_17) begin
                                    busy_bit_7 <= _GEN_23;
                                  end else if (_T_19) begin
                                    busy_bit_7 <= _GEN_23;
                                  end else if (_T_21) begin
                                    busy_bit_7 <= _GEN_39;
                                  end
                                end else if (_T_24) begin
                                  if (3'h7 == io_release_0_rd_addr) begin
                                    busy_bit_7 <= 1'h0;
                                  end else begin
                                    busy_bit_7 <= _GEN_63;
                                  end
                                end else if (_T_26) begin
                                  busy_bit_7 <= _GEN_87;
                                end else begin
                                  busy_bit_7 <= _GEN_63;
                                end
                              end else if (_T_31) begin
                                busy_bit_7 <= _GEN_135;
                              end else if (_T_17) begin
                                busy_bit_7 <= _GEN_71;
                              end else if (_T_24) begin
                                busy_bit_7 <= _GEN_71;
                              end else if (_T_26) begin
                                busy_bit_7 <= _GEN_87;
                              end else begin
                                busy_bit_7 <= _GEN_63;
                              end
                            end else if (_T_34) begin
                              if (3'h7 == io_release_0_rd_addr) begin
                                busy_bit_7 <= 1'h0;
                              end else if (_T_17) begin
                                if (3'h7 == io_release_0_rd_addr) begin
                                  busy_bit_7 <= 1'h0;
                                end else if (_T_17) begin
                                  busy_bit_7 <= _GEN_71;
                                end else if (_T_24) begin
                                  busy_bit_7 <= _GEN_71;
                                end else if (_T_26) begin
                                  busy_bit_7 <= _GEN_87;
                                end else begin
                                  busy_bit_7 <= _GEN_63;
                                end
                              end else if (_T_29) begin
                                if (3'h7 == io_release_0_rd_addr) begin
                                  busy_bit_7 <= 1'h0;
                                end else begin
                                  busy_bit_7 <= _GEN_111;
                                end
                              end else if (_T_31) begin
                                busy_bit_7 <= _GEN_135;
                              end else begin
                                busy_bit_7 <= _GEN_111;
                              end
                            end else if (_T_36) begin
                              busy_bit_7 <= _GEN_183;
                            end else if (_T_17) begin
                              busy_bit_7 <= _GEN_119;
                            end else if (_T_29) begin
                              busy_bit_7 <= _GEN_119;
                            end else if (_T_31) begin
                              busy_bit_7 <= _GEN_135;
                            end else begin
                              busy_bit_7 <= _GEN_111;
                            end
                          end else if (_T_39) begin
                            if (3'h7 == io_release_0_rd_addr) begin
                              busy_bit_7 <= 1'h0;
                            end else if (_T_17) begin
                              if (3'h7 == io_release_0_rd_addr) begin
                                busy_bit_7 <= 1'h0;
                              end else if (_T_17) begin
                                busy_bit_7 <= _GEN_119;
                              end else if (_T_29) begin
                                busy_bit_7 <= _GEN_119;
                              end else if (_T_31) begin
                                busy_bit_7 <= _GEN_135;
                              end else begin
                                busy_bit_7 <= _GEN_111;
                              end
                            end else if (_T_34) begin
                              if (3'h7 == io_release_0_rd_addr) begin
                                busy_bit_7 <= 1'h0;
                              end else begin
                                busy_bit_7 <= _GEN_159;
                              end
                            end else if (_T_36) begin
                              busy_bit_7 <= _GEN_183;
                            end else begin
                              busy_bit_7 <= _GEN_159;
                            end
                          end else if (_T_41) begin
                            busy_bit_7 <= _GEN_231;
                          end else if (_T_17) begin
                            busy_bit_7 <= _GEN_167;
                          end else if (_T_34) begin
                            busy_bit_7 <= _GEN_167;
                          end else if (_T_36) begin
                            busy_bit_7 <= _GEN_183;
                          end else begin
                            busy_bit_7 <= _GEN_159;
                          end
                        end else if (_T_44) begin
                          if (3'h7 == io_release_0_rd_addr) begin
                            busy_bit_7 <= 1'h0;
                          end else if (_T_17) begin
                            if (3'h7 == io_release_0_rd_addr) begin
                              busy_bit_7 <= 1'h0;
                            end else if (_T_17) begin
                              busy_bit_7 <= _GEN_167;
                            end else if (_T_34) begin
                              busy_bit_7 <= _GEN_167;
                            end else if (_T_36) begin
                              busy_bit_7 <= _GEN_183;
                            end else begin
                              busy_bit_7 <= _GEN_159;
                            end
                          end else if (_T_39) begin
                            if (3'h7 == io_release_0_rd_addr) begin
                              busy_bit_7 <= 1'h0;
                            end else begin
                              busy_bit_7 <= _GEN_207;
                            end
                          end else if (_T_41) begin
                            busy_bit_7 <= _GEN_231;
                          end else begin
                            busy_bit_7 <= _GEN_207;
                          end
                        end else if (_T_46) begin
                          busy_bit_7 <= _GEN_279;
                        end else if (_T_17) begin
                          busy_bit_7 <= _GEN_215;
                        end else if (_T_39) begin
                          busy_bit_7 <= _GEN_215;
                        end else if (_T_41) begin
                          busy_bit_7 <= _GEN_231;
                        end else begin
                          busy_bit_7 <= _GEN_207;
                        end
                      end else if (_T_49) begin
                        if (3'h7 == io_release_0_rd_addr) begin
                          busy_bit_7 <= 1'h0;
                        end else if (_T_17) begin
                          if (3'h7 == io_release_0_rd_addr) begin
                            busy_bit_7 <= 1'h0;
                          end else if (_T_17) begin
                            busy_bit_7 <= _GEN_215;
                          end else if (_T_39) begin
                            busy_bit_7 <= _GEN_215;
                          end else if (_T_41) begin
                            busy_bit_7 <= _GEN_231;
                          end else begin
                            busy_bit_7 <= _GEN_207;
                          end
                        end else if (_T_44) begin
                          if (3'h7 == io_release_0_rd_addr) begin
                            busy_bit_7 <= 1'h0;
                          end else begin
                            busy_bit_7 <= _GEN_255;
                          end
                        end else if (_T_46) begin
                          busy_bit_7 <= _GEN_279;
                        end else begin
                          busy_bit_7 <= _GEN_255;
                        end
                      end else if (_T_51) begin
                        busy_bit_7 <= _GEN_327;
                      end else if (_T_17) begin
                        busy_bit_7 <= _GEN_263;
                      end else if (_T_44) begin
                        busy_bit_7 <= _GEN_263;
                      end else if (_T_46) begin
                        busy_bit_7 <= _GEN_279;
                      end else begin
                        busy_bit_7 <= _GEN_255;
                      end
                    end else if (_T_54) begin
                      if (3'h7 == io_release_0_rd_addr) begin
                        busy_bit_7 <= 1'h0;
                      end else if (_T_17) begin
                        if (3'h7 == io_release_0_rd_addr) begin
                          busy_bit_7 <= 1'h0;
                        end else if (_T_17) begin
                          busy_bit_7 <= _GEN_263;
                        end else if (_T_44) begin
                          busy_bit_7 <= _GEN_263;
                        end else if (_T_46) begin
                          busy_bit_7 <= _GEN_279;
                        end else begin
                          busy_bit_7 <= _GEN_255;
                        end
                      end else if (_T_49) begin
                        if (3'h7 == io_release_0_rd_addr) begin
                          busy_bit_7 <= 1'h0;
                        end else begin
                          busy_bit_7 <= _GEN_303;
                        end
                      end else if (_T_51) begin
                        busy_bit_7 <= _GEN_327;
                      end else begin
                        busy_bit_7 <= _GEN_303;
                      end
                    end else if (_T_56) begin
                      busy_bit_7 <= _GEN_375;
                    end else if (_T_17) begin
                      busy_bit_7 <= _GEN_311;
                    end else if (_T_49) begin
                      busy_bit_7 <= _GEN_311;
                    end else if (_T_51) begin
                      busy_bit_7 <= _GEN_327;
                    end else begin
                      busy_bit_7 <= _GEN_303;
                    end
                  end else if (_T_21) begin
                    busy_bit_7 <= _GEN_423;
                  end else if (_T_17) begin
                    if (3'h7 == io_release_0_rd_addr) begin
                      busy_bit_7 <= 1'h0;
                    end else if (_T_17) begin
                      busy_bit_7 <= _GEN_311;
                    end else if (_T_49) begin
                      busy_bit_7 <= _GEN_311;
                    end else if (_T_51) begin
                      busy_bit_7 <= _GEN_327;
                    end else begin
                      busy_bit_7 <= _GEN_303;
                    end
                  end else if (_T_54) begin
                    if (3'h7 == io_release_0_rd_addr) begin
                      busy_bit_7 <= 1'h0;
                    end else begin
                      busy_bit_7 <= _GEN_351;
                    end
                  end else if (_T_56) begin
                    busy_bit_7 <= _GEN_375;
                  end else begin
                    busy_bit_7 <= _GEN_351;
                  end
                end else if (_T_26) begin
                  busy_bit_7 <= _GEN_471;
                end else if (_T_17) begin
                  if (_T_17) begin
                    busy_bit_7 <= _GEN_359;
                  end else if (_T_54) begin
                    busy_bit_7 <= _GEN_359;
                  end else if (_T_56) begin
                    busy_bit_7 <= _GEN_375;
                  end else begin
                    busy_bit_7 <= _GEN_351;
                  end
                end else if (_T_21) begin
                  busy_bit_7 <= _GEN_423;
                end else if (_T_17) begin
                  busy_bit_7 <= _GEN_359;
                end else if (_T_54) begin
                  busy_bit_7 <= _GEN_359;
                end else if (_T_56) begin
                  busy_bit_7 <= _GEN_375;
                end else begin
                  busy_bit_7 <= _GEN_351;
                end
              end else if (_T_31) begin
                busy_bit_7 <= _GEN_519;
              end else if (_T_17) begin
                if (_T_17) begin
                  busy_bit_7 <= _GEN_399;
                end else if (_T_21) begin
                  busy_bit_7 <= _GEN_423;
                end else begin
                  busy_bit_7 <= _GEN_399;
                end
              end else if (_T_26) begin
                busy_bit_7 <= _GEN_471;
              end else if (_T_17) begin
                busy_bit_7 <= _GEN_399;
              end else if (_T_21) begin
                busy_bit_7 <= _GEN_423;
              end else begin
                busy_bit_7 <= _GEN_399;
              end
            end else if (_T_36) begin
              busy_bit_7 <= _GEN_567;
            end else if (_T_17) begin
              if (_T_17) begin
                busy_bit_7 <= _GEN_447;
              end else if (_T_26) begin
                busy_bit_7 <= _GEN_471;
              end else begin
                busy_bit_7 <= _GEN_447;
              end
            end else if (_T_31) begin
              busy_bit_7 <= _GEN_519;
            end else if (_T_17) begin
              busy_bit_7 <= _GEN_447;
            end else if (_T_26) begin
              busy_bit_7 <= _GEN_471;
            end else begin
              busy_bit_7 <= _GEN_447;
            end
          end else if (_T_41) begin
            busy_bit_7 <= _GEN_615;
          end else if (_T_17) begin
            if (_T_17) begin
              busy_bit_7 <= _GEN_495;
            end else if (_T_31) begin
              busy_bit_7 <= _GEN_519;
            end else begin
              busy_bit_7 <= _GEN_495;
            end
          end else if (_T_36) begin
            busy_bit_7 <= _GEN_567;
          end else if (_T_17) begin
            busy_bit_7 <= _GEN_495;
          end else if (_T_31) begin
            busy_bit_7 <= _GEN_519;
          end else begin
            busy_bit_7 <= _GEN_495;
          end
        end else if (_T_46) begin
          busy_bit_7 <= _GEN_663;
        end else if (_T_17) begin
          if (_T_17) begin
            busy_bit_7 <= _GEN_543;
          end else if (_T_36) begin
            busy_bit_7 <= _GEN_567;
          end else begin
            busy_bit_7 <= _GEN_543;
          end
        end else if (_T_41) begin
          busy_bit_7 <= _GEN_615;
        end else if (_T_17) begin
          busy_bit_7 <= _GEN_543;
        end else if (_T_36) begin
          busy_bit_7 <= _GEN_567;
        end else begin
          busy_bit_7 <= _GEN_543;
        end
      end else if (_T_51) begin
        busy_bit_7 <= _GEN_711;
      end else if (_T_17) begin
        if (_T_17) begin
          busy_bit_7 <= _GEN_591;
        end else if (_T_41) begin
          busy_bit_7 <= _GEN_615;
        end else begin
          busy_bit_7 <= _GEN_591;
        end
      end else if (_T_46) begin
        busy_bit_7 <= _GEN_663;
      end else if (_T_17) begin
        busy_bit_7 <= _GEN_591;
      end else if (_T_41) begin
        busy_bit_7 <= _GEN_615;
      end else begin
        busy_bit_7 <= _GEN_591;
      end
    end else if (_T_56) begin
      busy_bit_7 <= _GEN_759;
    end else if (_T_17) begin
      if (_T_17) begin
        busy_bit_7 <= _GEN_639;
      end else if (_T_46) begin
        busy_bit_7 <= _GEN_663;
      end else begin
        busy_bit_7 <= _GEN_639;
      end
    end else if (_T_51) begin
      busy_bit_7 <= _GEN_711;
    end else if (_T_17) begin
      busy_bit_7 <= _GEN_639;
    end else if (_T_46) begin
      busy_bit_7 <= _GEN_663;
    end else begin
      busy_bit_7 <= _GEN_639;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"busy_bit: "); // @[BusyBit.scala 40:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",1'h0); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_1); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_2); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_3); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_4); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_5); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_6); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"%d, ",busy_bit_7); // @[BusyBit.scala 40:57]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_98) begin
          $fwrite(32'h80000002,"\n"); // @[BusyBit.scala 40:86]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ID(
  input         clock,
  input         reset,
  input         io_predict,
  input         io_branch_mispredicted,
  input         io_branch_graduated,
  input  [15:0] io_if_out_pc,
  input  [3:0]  io_if_out_inst_bits_op,
  input  [2:0]  io_if_out_inst_bits_rd,
  input  [2:0]  io_if_out_inst_bits_rs,
  input  [5:0]  io_if_out_inst_bits_disp6u,
  input  [2:0]  io_commit_0_rd_addr,
  input         io_commit_0_rf_w,
  input  [15:0] io_commit_0_data,
  input         io_unreserved_head_0_valid,
  input  [3:0]  io_unreserved_head_0_bits,
  output        io_used_num,
  output [15:0] io_jump_pc,
  output [15:0] io_next_pc,
  output        io_inst_info_valid,
  output [2:0]  io_inst_info_rd_addr,
  output [3:0]  io_inst_info_rob_addr,
  output [2:0]  io_inst_info_ctrl_alu_op,
  output        io_inst_info_ctrl_is_jump,
  output        io_inst_info_ctrl_is_branch,
  output        io_inst_info_ctrl_rf_w,
  output        io_inst_info_ctrl_mem_r,
  output        io_inst_info_ctrl_mem_w,
  output [15:0] io_source_0,
  output [15:0] io_source_1,
  output [15:0] io_rd,
  output        io_stall,
  output [15:0] io_pc,
  output [15:0] io_rf4debug_1,
  output [15:0] io_rf4debug_2,
  output [15:0] io_rf4debug_3,
  output [15:0] io_rf4debug_4,
  output [15:0] io_rf4debug_5,
  output [15:0] io_rf4debug_6,
  output [15:0] io_rf4debug_7
);
  wire [3:0] decoder_io_inst_bits_op; // @[ID.scala 49:32]
  wire [2:0] decoder_io_ctrl_alu_op; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_is_jump; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_is_branch; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_rf_w; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_mem_r; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_mem_w; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_rs1_use; // @[ID.scala 49:32]
  wire  decoder_io_ctrl_rs2_use; // @[ID.scala 49:32]
  wire [15:0] decoder_io_source_sel_0; // @[ID.scala 49:32]
  wire [15:0] decoder_io_source_sel_1; // @[ID.scala 49:32]
  wire  reg_file_clock; // @[ID.scala 52:38]
  wire  reg_file_reset; // @[ID.scala 52:38]
  wire [2:0] reg_file_io_read_addr_0; // @[ID.scala 52:38]
  wire [2:0] reg_file_io_read_addr_1; // @[ID.scala 52:38]
  wire [2:0] reg_file_io_write_0_rd_addr; // @[ID.scala 52:38]
  wire  reg_file_io_write_0_rf_w; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_write_0_data; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_out_0; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_out_1; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_1; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_2; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_3; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_4; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_5; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_6; // @[ID.scala 52:38]
  wire [15:0] reg_file_io_rf4debug_7; // @[ID.scala 52:38]
  wire  busy_bit_clock; // @[ID.scala 57:33]
  wire  busy_bit_reset; // @[ID.scala 57:33]
  wire  busy_bit_io_branch_mispredicted; // @[ID.scala 57:33]
  wire  busy_bit_io_branch_graduated; // @[ID.scala 57:33]
  wire [2:0] busy_bit_io_release_0_rd_addr; // @[ID.scala 57:33]
  wire  busy_bit_io_release_0_rf_w; // @[ID.scala 57:33]
  wire [2:0] busy_bit_io_req_rs_addr_0; // @[ID.scala 57:33]
  wire [2:0] busy_bit_io_req_rs_addr_1; // @[ID.scala 57:33]
  wire  busy_bit_io_req_rd_w; // @[ID.scala 57:33]
  wire [2:0] busy_bit_io_req_rd_addr; // @[ID.scala 57:33]
  wire  busy_bit_io_rs_available_0; // @[ID.scala 57:33]
  wire  busy_bit_io_rs_available_1; // @[ID.scala 57:33]
  reg [15:0] if_out_r_pc; // @[ID.scala 37:32]
  reg [31:0] _RAND_0;
  reg [3:0] if_out_r_inst_bits_op; // @[ID.scala 37:32]
  reg [31:0] _RAND_1;
  reg [2:0] if_out_r_inst_bits_rd; // @[ID.scala 37:32]
  reg [31:0] _RAND_2;
  reg [2:0] if_out_r_inst_bits_rs; // @[ID.scala 37:32]
  reg [31:0] _RAND_3;
  reg [5:0] if_out_r_inst_bits_disp6u; // @[ID.scala 37:32]
  reg [31:0] _RAND_4;
  wire [15:0] if_out_pc; // @[ID.scala 38:16]
  wire [3:0] if_out_inst_bits_op; // @[ID.scala 38:16]
  wire [2:0] if_out_inst_bits_rs; // @[ID.scala 38:16]
  wire [5:0] if_out_inst_bits_disp6u; // @[ID.scala 38:16]
  reg  predict_r; // @[ID.scala 41:32]
  reg [31:0] _RAND_5;
  wire  predict; // @[ID.scala 42:17]
  reg  _T_8; // @[ID.scala 75:16]
  reg [31:0] _RAND_6;
  wire  _T_9; // @[ID.scala 75:5]
  reg  _T_12; // @[ID.scala 76:16]
  reg [31:0] _RAND_7;
  wire  _T_13; // @[ID.scala 76:75]
  wire  clear_instruction; // @[ID.scala 76:5]
  wire  _T_2; // @[ID.scala 65:27]
  wire  _T_15; // @[ID.scala 85:37]
  wire  _T_16; // @[ID.scala 85:34]
  wire  _T_17; // @[ID.scala 86:37]
  wire  _T_18; // @[ID.scala 86:34]
  wire  operands_available; // @[ID.scala 85:63]
  wire  _T_19; // @[ID.scala 96:44]
  wire  _T_20; // @[ID.scala 96:67]
  wire  _T_21; // @[ID.scala 96:64]
  wire  stall; // @[ID.scala 96:15]
  wire  _T_3; // @[ID.scala 65:49]
  wire  _T_4; // @[ID.scala 65:46]
  wire  _T_7; // @[ID.scala 75:36]
  wire  _T_11; // @[ID.scala 76:36]
  reg  _T_23; // @[ID.scala 97:22]
  reg [31:0] _RAND_8;
  wire  _T_24; // @[ID.scala 101:11]
  wire  _T_25; // @[ID.scala 101:55]
  wire  _T_26; // @[ID.scala 101:32]
  reg  _T_28; // @[ID.scala 100:25]
  reg [31:0] _RAND_9;
  wire  _T_32; // @[ID.scala 107:5]
  reg  _T_35; // @[ID.scala 106:32]
  reg [31:0] _RAND_10;
  reg [2:0] _T_44; // @[ID.scala 112:34]
  reg [31:0] _RAND_11;
  reg [2:0] _T_51_alu_op; // @[ID.scala 114:31]
  reg [31:0] _RAND_12;
  reg  _T_51_is_jump; // @[ID.scala 114:31]
  reg [31:0] _RAND_13;
  reg  _T_51_is_branch; // @[ID.scala 114:31]
  reg [31:0] _RAND_14;
  reg  _T_51_rf_w; // @[ID.scala 114:31]
  reg [31:0] _RAND_15;
  reg  _T_51_mem_r; // @[ID.scala 114:31]
  reg [31:0] _RAND_16;
  reg  _T_51_mem_w; // @[ID.scala 114:31]
  reg [31:0] _RAND_17;
  wire [8:0] _T_52; // @[Cat.scala 29:58]
  wire  _T_56; // @[InstBits.scala 18:43]
  wire [6:0] _T_57; // @[InstBits.scala 18:28]
  wire [15:0] _T_59; // @[Cat.scala 29:58]
  wire [15:0] _T_61; // @[ID.scala 120:15]
  wire  _T_65; // @[InstBits.scala 16:45]
  wire [9:0] _T_66; // @[InstBits.scala 16:29]
  wire [15:0] _T_67; // @[Cat.scala 29:58]
  wire [15:0] _T_69; // @[ID.scala 120:51]
  reg [15:0] _T_71; // @[ID.scala 119:24]
  reg [31:0] _RAND_18;
  reg [15:0] _T_74; // @[ID.scala 122:24]
  reg [31:0] _RAND_19;
  wire  _T_77; // @[Mux.scala 68:19]
  wire  _T_79; // @[Mux.scala 68:19]
  reg [15:0] _T_81; // @[ID.scala 124:26]
  reg [31:0] _RAND_20;
  wire  _T_90; // @[Mux.scala 68:19]
  wire  _T_92; // @[Mux.scala 68:19]
  wire  _T_94; // @[Mux.scala 68:19]
  reg [15:0] _T_96; // @[ID.scala 129:26]
  reg [31:0] _RAND_21;
  reg [15:0] _T_97; // @[ID.scala 134:19]
  reg [31:0] _RAND_22;
  reg [15:0] _T_98; // @[ID.scala 135:19]
  reg [31:0] _RAND_23;
  wire  _T_99; // @[ID.scala 137:9]
  wire  _T_100; // @[ID.scala 137:9]
  Decoder decoder ( // @[ID.scala 49:32]
    .io_inst_bits_op(decoder_io_inst_bits_op),
    .io_ctrl_alu_op(decoder_io_ctrl_alu_op),
    .io_ctrl_is_jump(decoder_io_ctrl_is_jump),
    .io_ctrl_is_branch(decoder_io_ctrl_is_branch),
    .io_ctrl_rf_w(decoder_io_ctrl_rf_w),
    .io_ctrl_mem_r(decoder_io_ctrl_mem_r),
    .io_ctrl_mem_w(decoder_io_ctrl_mem_w),
    .io_ctrl_rs1_use(decoder_io_ctrl_rs1_use),
    .io_ctrl_rs2_use(decoder_io_ctrl_rs2_use),
    .io_source_sel_0(decoder_io_source_sel_0),
    .io_source_sel_1(decoder_io_source_sel_1)
  );
  RegisterFile reg_file ( // @[ID.scala 52:38]
    .clock(reg_file_clock),
    .reset(reg_file_reset),
    .io_read_addr_0(reg_file_io_read_addr_0),
    .io_read_addr_1(reg_file_io_read_addr_1),
    .io_write_0_rd_addr(reg_file_io_write_0_rd_addr),
    .io_write_0_rf_w(reg_file_io_write_0_rf_w),
    .io_write_0_data(reg_file_io_write_0_data),
    .io_out_0(reg_file_io_out_0),
    .io_out_1(reg_file_io_out_1),
    .io_rf4debug_1(reg_file_io_rf4debug_1),
    .io_rf4debug_2(reg_file_io_rf4debug_2),
    .io_rf4debug_3(reg_file_io_rf4debug_3),
    .io_rf4debug_4(reg_file_io_rf4debug_4),
    .io_rf4debug_5(reg_file_io_rf4debug_5),
    .io_rf4debug_6(reg_file_io_rf4debug_6),
    .io_rf4debug_7(reg_file_io_rf4debug_7)
  );
  BusyBit busy_bit ( // @[ID.scala 57:33]
    .clock(busy_bit_clock),
    .reset(busy_bit_reset),
    .io_branch_mispredicted(busy_bit_io_branch_mispredicted),
    .io_branch_graduated(busy_bit_io_branch_graduated),
    .io_release_0_rd_addr(busy_bit_io_release_0_rd_addr),
    .io_release_0_rf_w(busy_bit_io_release_0_rf_w),
    .io_req_rs_addr_0(busy_bit_io_req_rs_addr_0),
    .io_req_rs_addr_1(busy_bit_io_req_rs_addr_1),
    .io_req_rd_w(busy_bit_io_req_rd_w),
    .io_req_rd_addr(busy_bit_io_req_rd_addr),
    .io_rs_available_0(busy_bit_io_rs_available_0),
    .io_rs_available_1(busy_bit_io_rs_available_1)
  );
  assign if_out_pc = io_stall ? if_out_r_pc : io_if_out_pc; // @[ID.scala 38:16]
  assign if_out_inst_bits_op = io_stall ? if_out_r_inst_bits_op : io_if_out_inst_bits_op; // @[ID.scala 38:16]
  assign if_out_inst_bits_rs = io_stall ? if_out_r_inst_bits_rs : io_if_out_inst_bits_rs; // @[ID.scala 38:16]
  assign if_out_inst_bits_disp6u = io_stall ? if_out_r_inst_bits_disp6u : io_if_out_inst_bits_disp6u; // @[ID.scala 38:16]
  assign predict = io_stall ? predict_r : io_predict; // @[ID.scala 42:17]
  assign _T_9 = io_branch_mispredicted | _T_8; // @[ID.scala 75:5]
  assign _T_13 = _T_12 & predict; // @[ID.scala 76:75]
  assign clear_instruction = _T_9 | _T_13; // @[ID.scala 76:5]
  assign _T_2 = clear_instruction == 1'h0; // @[ID.scala 65:27]
  assign _T_15 = decoder_io_ctrl_rs1_use == 1'h0; // @[ID.scala 85:37]
  assign _T_16 = busy_bit_io_rs_available_0 | _T_15; // @[ID.scala 85:34]
  assign _T_17 = decoder_io_ctrl_rs2_use == 1'h0; // @[ID.scala 86:37]
  assign _T_18 = busy_bit_io_rs_available_1 | _T_17; // @[ID.scala 86:34]
  assign operands_available = _T_16 & _T_18; // @[ID.scala 85:63]
  assign _T_19 = operands_available == 1'h0; // @[ID.scala 96:44]
  assign _T_20 = io_unreserved_head_0_valid == 1'h0; // @[ID.scala 96:67]
  assign _T_21 = _T_19 | _T_20; // @[ID.scala 96:64]
  assign stall = clear_instruction ? 1'h0 : _T_21; // @[ID.scala 96:15]
  assign _T_3 = stall == 1'h0; // @[ID.scala 65:49]
  assign _T_4 = _T_2 & _T_3; // @[ID.scala 65:46]
  assign _T_7 = _T_2 & decoder_io_ctrl_is_jump; // @[ID.scala 75:36]
  assign _T_11 = _T_2 & decoder_io_ctrl_is_branch; // @[ID.scala 76:36]
  assign _T_24 = stall | clear_instruction; // @[ID.scala 101:11]
  assign _T_25 = if_out_inst_bits_op == 4'h0; // @[ID.scala 101:55]
  assign _T_26 = _T_24 | _T_25; // @[ID.scala 101:32]
  assign _T_32 = _T_26 == 1'h0; // @[ID.scala 107:5]
  assign _T_52 = {if_out_inst_bits_rs,if_out_inst_bits_disp6u}; // @[Cat.scala 29:58]
  assign _T_56 = _T_52[8]; // @[InstBits.scala 18:43]
  assign _T_57 = _T_56 ? 7'h7f : 7'h0; // @[InstBits.scala 18:28]
  assign _T_59 = {_T_57,if_out_inst_bits_rs,if_out_inst_bits_disp6u}; // @[Cat.scala 29:58]
  assign _T_61 = if_out_pc + _T_59; // @[ID.scala 120:15]
  assign _T_65 = if_out_inst_bits_disp6u[5]; // @[InstBits.scala 16:45]
  assign _T_66 = _T_65 ? 10'h3ff : 10'h0; // @[InstBits.scala 16:29]
  assign _T_67 = {_T_66,if_out_inst_bits_disp6u}; // @[Cat.scala 29:58]
  assign _T_69 = if_out_pc + _T_67; // @[ID.scala 120:51]
  assign _T_77 = 16'h1 == decoder_io_source_sel_0; // @[Mux.scala 68:19]
  assign _T_79 = 16'h3 == decoder_io_source_sel_0; // @[Mux.scala 68:19]
  assign _T_90 = 16'h0 == decoder_io_source_sel_1; // @[Mux.scala 68:19]
  assign _T_92 = 16'h1 == decoder_io_source_sel_1; // @[Mux.scala 68:19]
  assign _T_94 = 16'h2 == decoder_io_source_sel_1; // @[Mux.scala 68:19]
  assign _T_99 = $unsigned(reset); // @[ID.scala 137:9]
  assign _T_100 = _T_99 == 1'h0; // @[ID.scala 137:9]
  assign io_used_num = _T_28; // @[ID.scala 100:15]
  assign io_jump_pc = _T_71; // @[ID.scala 119:14]
  assign io_next_pc = _T_74; // @[ID.scala 122:14]
  assign io_inst_info_valid = _T_35; // @[ID.scala 106:22]
  assign io_inst_info_rd_addr = _T_44; // @[ID.scala 112:24]
  assign io_inst_info_rob_addr = io_unreserved_head_0_bits; // @[ID.scala 113:25]
  assign io_inst_info_ctrl_alu_op = _T_51_alu_op; // @[ID.scala 114:21]
  assign io_inst_info_ctrl_is_jump = _T_51_is_jump; // @[ID.scala 114:21]
  assign io_inst_info_ctrl_is_branch = _T_51_is_branch; // @[ID.scala 114:21]
  assign io_inst_info_ctrl_rf_w = _T_51_rf_w; // @[ID.scala 114:21]
  assign io_inst_info_ctrl_mem_r = _T_51_mem_r; // @[ID.scala 114:21]
  assign io_inst_info_ctrl_mem_w = _T_51_mem_w; // @[ID.scala 114:21]
  assign io_source_0 = _T_81; // @[ID.scala 124:16]
  assign io_source_1 = _T_96; // @[ID.scala 129:16]
  assign io_rd = _T_97; // @[ID.scala 134:9]
  assign io_stall = _T_23; // @[ID.scala 97:12]
  assign io_pc = _T_98; // @[ID.scala 135:9]
  assign io_rf4debug_1 = reg_file_io_rf4debug_1; // @[ID.scala 145:15]
  assign io_rf4debug_2 = reg_file_io_rf4debug_2; // @[ID.scala 145:15]
  assign io_rf4debug_3 = reg_file_io_rf4debug_3; // @[ID.scala 145:15]
  assign io_rf4debug_4 = reg_file_io_rf4debug_4; // @[ID.scala 145:15]
  assign io_rf4debug_5 = reg_file_io_rf4debug_5; // @[ID.scala 145:15]
  assign io_rf4debug_6 = reg_file_io_rf4debug_6; // @[ID.scala 145:15]
  assign io_rf4debug_7 = reg_file_io_rf4debug_7; // @[ID.scala 145:15]
  assign decoder_io_inst_bits_op = io_stall ? if_out_r_inst_bits_op : io_if_out_inst_bits_op; // @[ID.scala 50:24]
  assign reg_file_clock = clock;
  assign reg_file_reset = reset;
  assign reg_file_io_read_addr_0 = io_stall ? if_out_r_inst_bits_rd : io_if_out_inst_bits_rd; // @[ID.scala 53:28]
  assign reg_file_io_read_addr_1 = io_stall ? if_out_r_inst_bits_rs : io_if_out_inst_bits_rs; // @[ID.scala 54:28]
  assign reg_file_io_write_0_rd_addr = io_commit_0_rd_addr; // @[ID.scala 55:21]
  assign reg_file_io_write_0_rf_w = io_commit_0_rf_w; // @[ID.scala 55:21]
  assign reg_file_io_write_0_data = io_commit_0_data; // @[ID.scala 55:21]
  assign busy_bit_clock = clock;
  assign busy_bit_reset = reset;
  assign busy_bit_io_branch_mispredicted = io_branch_mispredicted; // @[ID.scala 58:35]
  assign busy_bit_io_branch_graduated = io_branch_graduated; // @[ID.scala 59:32]
  assign busy_bit_io_release_0_rd_addr = io_commit_0_rd_addr; // @[ID.scala 60:23]
  assign busy_bit_io_release_0_rf_w = io_commit_0_rf_w; // @[ID.scala 60:23]
  assign busy_bit_io_req_rs_addr_0 = io_stall ? if_out_r_inst_bits_rd : io_if_out_inst_bits_rd; // @[ID.scala 61:30]
  assign busy_bit_io_req_rs_addr_1 = io_stall ? if_out_r_inst_bits_rs : io_if_out_inst_bits_rs; // @[ID.scala 62:30]
  assign busy_bit_io_req_rd_w = _T_4 & decoder_io_ctrl_rf_w; // @[ID.scala 65:24]
  assign busy_bit_io_req_rd_addr = io_stall ? if_out_r_inst_bits_rd : io_if_out_inst_bits_rd; // @[ID.scala 66:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_out_r_pc = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  if_out_r_inst_bits_op = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  if_out_r_inst_bits_rd = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  if_out_r_inst_bits_rs = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  if_out_r_inst_bits_disp6u = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  predict_r = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_8 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_12 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_23 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_28 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_35 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_44 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_51_alu_op = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_51_is_jump = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_51_is_branch = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_51_rf_w = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_51_mem_r = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_51_mem_w = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_71 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_74 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_81 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_96 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_97 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_98 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (!(io_stall)) begin
      if_out_r_pc <= io_if_out_pc;
    end
    if (!(io_stall)) begin
      if_out_r_inst_bits_op <= io_if_out_inst_bits_op;
    end
    if (!(io_stall)) begin
      if_out_r_inst_bits_rd <= io_if_out_inst_bits_rd;
    end
    if (!(io_stall)) begin
      if_out_r_inst_bits_rs <= io_if_out_inst_bits_rs;
    end
    if (!(io_stall)) begin
      if_out_r_inst_bits_disp6u <= io_if_out_inst_bits_disp6u;
    end
    if (!(io_stall)) begin
      predict_r <= io_predict;
    end
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      _T_8 <= _T_7;
    end
    if (reset) begin
      _T_12 <= 1'h0;
    end else begin
      _T_12 <= _T_11;
    end
    if (reset) begin
      _T_23 <= 1'h0;
    end else if (clear_instruction) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else if (_T_26) begin
      _T_28 <= 1'h0;
    end else begin
      _T_28 <= 1'h1;
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      _T_35 <= _T_32;
    end
    if (reset) begin
      _T_44 <= 3'h0;
    end else if (io_stall) begin
      _T_44 <= if_out_r_inst_bits_rd;
    end else begin
      _T_44 <= io_if_out_inst_bits_rd;
    end
    if (reset) begin
      _T_51_alu_op <= 3'h0;
    end else if (_T_24) begin
      _T_51_alu_op <= 3'h0;
    end else begin
      _T_51_alu_op <= decoder_io_ctrl_alu_op;
    end
    if (reset) begin
      _T_51_is_jump <= 1'h0;
    end else if (_T_24) begin
      _T_51_is_jump <= 1'h0;
    end else begin
      _T_51_is_jump <= decoder_io_ctrl_is_jump;
    end
    if (reset) begin
      _T_51_is_branch <= 1'h0;
    end else if (_T_24) begin
      _T_51_is_branch <= 1'h0;
    end else begin
      _T_51_is_branch <= decoder_io_ctrl_is_branch;
    end
    if (reset) begin
      _T_51_rf_w <= 1'h0;
    end else if (_T_24) begin
      _T_51_rf_w <= 1'h0;
    end else begin
      _T_51_rf_w <= decoder_io_ctrl_rf_w;
    end
    if (reset) begin
      _T_51_mem_r <= 1'h0;
    end else if (_T_24) begin
      _T_51_mem_r <= 1'h0;
    end else begin
      _T_51_mem_r <= decoder_io_ctrl_mem_r;
    end
    if (reset) begin
      _T_51_mem_w <= 1'h0;
    end else if (_T_24) begin
      _T_51_mem_w <= 1'h0;
    end else begin
      _T_51_mem_w <= decoder_io_ctrl_mem_w;
    end
    if (decoder_io_ctrl_is_jump) begin
      _T_71 <= _T_61;
    end else begin
      _T_71 <= _T_69;
    end
    _T_74 <= if_out_pc + 16'h1;
    if (_T_79) begin
      _T_81 <= {{10'd0}, if_out_inst_bits_disp6u};
    end else if (_T_77) begin
      _T_81 <= reg_file_io_out_0;
    end else begin
      _T_81 <= 16'h0;
    end
    if (_T_94) begin
      _T_96 <= _T_59;
    end else if (_T_92) begin
      _T_96 <= reg_file_io_out_1;
    end else begin
      _T_96 <= {{15'd0}, _T_90};
    end
    _T_97 <= reg_file_io_out_0;
    if (io_stall) begin
      _T_98 <= if_out_r_pc;
    end else begin
      _T_98 <= io_if_out_pc;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"branch_mispredicted_enable: %d, branch_mispredicted: %d\n",io_branch_graduated,io_branch_mispredicted); // @[ID.scala 137:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"stall: %d, !operands_avail: %d, !rob_avail(0): %d\n",stall,_T_19,_T_20); // @[ID.scala 138:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"source(0): %d\n",io_source_0); // @[ID.scala 140:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"source(1): %d\n",io_source_1); // @[ID.scala 141:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"next_addr: %d\n",io_jump_pc); // @[ID.scala 142:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"----------\n"); // @[ID.scala 143:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_inst_info_valid,
  input  [2:0]  io_inst_info_rd_addr,
  input  [3:0]  io_inst_info_rob_addr,
  input  [2:0]  io_inst_info_ctrl_alu_op,
  input         io_inst_info_ctrl_is_branch,
  input         io_inst_info_ctrl_rf_w,
  input         io_inst_info_ctrl_mem_r,
  input         io_inst_info_ctrl_mem_w,
  input  [15:0] io_source_0,
  input  [15:0] io_source_1,
  input  [15:0] io_next_pc,
  input  [15:0] io_branch_pc,
  input  [15:0] io_rd,
  input         io_predict,
  input  [15:0] io_pc,
  output [15:0] io_alu_out,
  output        io_inst_info_out_valid,
  output [2:0]  io_inst_info_out_rd_addr,
  output [3:0]  io_inst_info_out_rob_addr,
  output        io_inst_info_out_ctrl_is_branch,
  output        io_inst_info_out_ctrl_rf_w,
  output        io_inst_info_out_ctrl_mem_r,
  output        io_inst_info_out_ctrl_mem_w,
  output [15:0] io_restoration_pc,
  output [15:0] io_rd_out,
  output [15:0] io_pc_out,
  output        io_mispredicted
);
  wire [15:0] _T_1; // @[ALU.scala 29:34]
  wire [15:0] _T_3; // @[ALU.scala 30:34]
  wire [15:0] _T_4; // @[ALU.scala 31:34]
  wire [15:0] _T_5; // @[ALU.scala 32:34]
  wire  _T_6; // @[ALU.scala 33:37]
  wire  _T_7; // @[ALU.scala 34:35]
  wire  _T_8; // @[Mux.scala 68:19]
  wire  _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire  _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [15:0] _T_13; // @[Mux.scala 68:16]
  wire  _T_14; // @[Mux.scala 68:19]
  wire [15:0] _T_15; // @[Mux.scala 68:16]
  wire  _T_16; // @[Mux.scala 68:19]
  wire [15:0] _T_17; // @[Mux.scala 68:16]
  wire  _T_18; // @[Mux.scala 68:19]
  wire [15:0] alu_out; // @[Mux.scala 68:16]
  reg [15:0] _T_19; // @[ALU.scala 36:24]
  reg [31:0] _RAND_0;
  reg  _T_22_valid; // @[ALU.scala 37:30]
  reg [31:0] _RAND_1;
  reg [2:0] _T_22_rd_addr; // @[ALU.scala 37:30]
  reg [31:0] _RAND_2;
  reg [3:0] _T_22_rob_addr; // @[ALU.scala 37:30]
  reg [31:0] _RAND_3;
  reg  _T_22_ctrl_is_branch; // @[ALU.scala 37:30]
  reg [31:0] _RAND_4;
  reg  _T_22_ctrl_rf_w; // @[ALU.scala 37:30]
  reg [31:0] _RAND_5;
  reg  _T_22_ctrl_mem_r; // @[ALU.scala 37:30]
  reg [31:0] _RAND_6;
  reg  _T_22_ctrl_mem_w; // @[ALU.scala 37:30]
  reg [31:0] _RAND_7;
  reg [15:0] _T_24; // @[ALU.scala 38:31]
  reg [31:0] _RAND_8;
  reg [15:0] _T_25; // @[ALU.scala 42:23]
  reg [31:0] _RAND_9;
  reg [15:0] _T_26; // @[ALU.scala 43:23]
  reg [31:0] _RAND_10;
  wire [15:0] _GEN_0; // @[ALU.scala 44:73]
  wire  _T_27; // @[ALU.scala 44:73]
  reg  _T_29; // @[ALU.scala 44:29]
  reg [31:0] _RAND_11;
  assign _T_1 = io_source_0 + io_source_1; // @[ALU.scala 29:34]
  assign _T_3 = io_source_0 - io_source_1; // @[ALU.scala 30:34]
  assign _T_4 = io_source_0 & io_source_1; // @[ALU.scala 31:34]
  assign _T_5 = io_source_0 | io_source_1; // @[ALU.scala 32:34]
  assign _T_6 = io_source_0 == io_source_1; // @[ALU.scala 33:37]
  assign _T_7 = io_source_0 > io_source_1; // @[ALU.scala 34:35]
  assign _T_8 = 3'h5 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 & _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h4 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? _T_6 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 3'h3 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign _T_13 = _T_12 ? _T_5 : {{15'd0}, _T_11}; // @[Mux.scala 68:16]
  assign _T_14 = 3'h2 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign _T_15 = _T_14 ? _T_4 : _T_13; // @[Mux.scala 68:16]
  assign _T_16 = 3'h1 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign _T_17 = _T_16 ? _T_3 : _T_15; // @[Mux.scala 68:16]
  assign _T_18 = 3'h0 == io_inst_info_ctrl_alu_op; // @[Mux.scala 68:19]
  assign alu_out = _T_18 ? _T_1 : _T_17; // @[Mux.scala 68:16]
  assign _GEN_0 = {{15'd0}, io_predict}; // @[ALU.scala 44:73]
  assign _T_27 = _GEN_0 != alu_out; // @[ALU.scala 44:73]
  assign io_alu_out = _T_19; // @[ALU.scala 36:14]
  assign io_inst_info_out_valid = _T_22_valid; // @[ALU.scala 37:20]
  assign io_inst_info_out_rd_addr = _T_22_rd_addr; // @[ALU.scala 37:20]
  assign io_inst_info_out_rob_addr = _T_22_rob_addr; // @[ALU.scala 37:20]
  assign io_inst_info_out_ctrl_is_branch = _T_22_ctrl_is_branch; // @[ALU.scala 37:20]
  assign io_inst_info_out_ctrl_rf_w = _T_22_ctrl_rf_w; // @[ALU.scala 37:20]
  assign io_inst_info_out_ctrl_mem_r = _T_22_ctrl_mem_r; // @[ALU.scala 37:20]
  assign io_inst_info_out_ctrl_mem_w = _T_22_ctrl_mem_w; // @[ALU.scala 37:20]
  assign io_restoration_pc = _T_24; // @[ALU.scala 38:21]
  assign io_rd_out = _T_25; // @[ALU.scala 42:13]
  assign io_pc_out = _T_26; // @[ALU.scala 43:13]
  assign io_mispredicted = _T_29; // @[ALU.scala 44:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_22_rd_addr = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_22_rob_addr = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_22_ctrl_is_branch = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_22_ctrl_rf_w = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22_ctrl_mem_r = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_22_ctrl_mem_w = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_24 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_25 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_26 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_29 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_18) begin
      _T_19 <= _T_1;
    end else if (_T_16) begin
      _T_19 <= _T_3;
    end else if (_T_14) begin
      _T_19 <= _T_4;
    end else if (_T_12) begin
      _T_19 <= _T_5;
    end else begin
      _T_19 <= {{15'd0}, _T_11};
    end
    if (reset) begin
      _T_22_valid <= 1'h0;
    end else begin
      _T_22_valid <= io_inst_info_valid;
    end
    if (reset) begin
      _T_22_rd_addr <= 3'h0;
    end else begin
      _T_22_rd_addr <= io_inst_info_rd_addr;
    end
    if (reset) begin
      _T_22_rob_addr <= 4'h0;
    end else begin
      _T_22_rob_addr <= io_inst_info_rob_addr;
    end
    if (reset) begin
      _T_22_ctrl_is_branch <= 1'h0;
    end else begin
      _T_22_ctrl_is_branch <= io_inst_info_ctrl_is_branch;
    end
    if (reset) begin
      _T_22_ctrl_rf_w <= 1'h0;
    end else begin
      _T_22_ctrl_rf_w <= io_inst_info_ctrl_rf_w;
    end
    if (reset) begin
      _T_22_ctrl_mem_r <= 1'h0;
    end else begin
      _T_22_ctrl_mem_r <= io_inst_info_ctrl_mem_r;
    end
    if (reset) begin
      _T_22_ctrl_mem_w <= 1'h0;
    end else begin
      _T_22_ctrl_mem_w <= io_inst_info_ctrl_mem_w;
    end
    if (io_predict) begin
      _T_24 <= io_next_pc;
    end else begin
      _T_24 <= io_branch_pc;
    end
    _T_25 <= io_rd;
    _T_26 <= io_pc;
    _T_29 <= io_inst_info_ctrl_is_branch & _T_27;
  end
endmodule
module EX(
  input         clock,
  input         reset,
  input         io_inst_info_valid,
  input  [2:0]  io_inst_info_rd_addr,
  input  [3:0]  io_inst_info_rob_addr,
  input  [2:0]  io_inst_info_ctrl_alu_op,
  input         io_inst_info_ctrl_is_branch,
  input         io_inst_info_ctrl_rf_w,
  input         io_inst_info_ctrl_mem_r,
  input         io_inst_info_ctrl_mem_w,
  input  [15:0] io_source_0,
  input  [15:0] io_source_1,
  input  [15:0] io_branch_pc,
  input  [15:0] io_next_pc,
  input  [15:0] io_rd,
  input         io_predict,
  input  [15:0] io_pc,
  output [15:0] io_alu_out,
  output        io_inst_info_out_valid,
  output [2:0]  io_inst_info_out_rd_addr,
  output [3:0]  io_inst_info_out_rob_addr,
  output        io_inst_info_out_ctrl_is_branch,
  output        io_inst_info_out_ctrl_rf_w,
  output        io_inst_info_out_ctrl_mem_r,
  output        io_inst_info_out_ctrl_mem_w,
  output [15:0] io_restoration_pc_out,
  output [15:0] io_rd_out,
  output [15:0] io_pc_out,
  output        io_mispredicted
);
  wire  alu_clock; // @[EX.scala 30:24]
  wire  alu_reset; // @[EX.scala 30:24]
  wire  alu_io_inst_info_valid; // @[EX.scala 30:24]
  wire [2:0] alu_io_inst_info_rd_addr; // @[EX.scala 30:24]
  wire [3:0] alu_io_inst_info_rob_addr; // @[EX.scala 30:24]
  wire [2:0] alu_io_inst_info_ctrl_alu_op; // @[EX.scala 30:24]
  wire  alu_io_inst_info_ctrl_is_branch; // @[EX.scala 30:24]
  wire  alu_io_inst_info_ctrl_rf_w; // @[EX.scala 30:24]
  wire  alu_io_inst_info_ctrl_mem_r; // @[EX.scala 30:24]
  wire  alu_io_inst_info_ctrl_mem_w; // @[EX.scala 30:24]
  wire [15:0] alu_io_source_0; // @[EX.scala 30:24]
  wire [15:0] alu_io_source_1; // @[EX.scala 30:24]
  wire [15:0] alu_io_next_pc; // @[EX.scala 30:24]
  wire [15:0] alu_io_branch_pc; // @[EX.scala 30:24]
  wire [15:0] alu_io_rd; // @[EX.scala 30:24]
  wire  alu_io_predict; // @[EX.scala 30:24]
  wire [15:0] alu_io_pc; // @[EX.scala 30:24]
  wire [15:0] alu_io_alu_out; // @[EX.scala 30:24]
  wire  alu_io_inst_info_out_valid; // @[EX.scala 30:24]
  wire [2:0] alu_io_inst_info_out_rd_addr; // @[EX.scala 30:24]
  wire [3:0] alu_io_inst_info_out_rob_addr; // @[EX.scala 30:24]
  wire  alu_io_inst_info_out_ctrl_is_branch; // @[EX.scala 30:24]
  wire  alu_io_inst_info_out_ctrl_rf_w; // @[EX.scala 30:24]
  wire  alu_io_inst_info_out_ctrl_mem_r; // @[EX.scala 30:24]
  wire  alu_io_inst_info_out_ctrl_mem_w; // @[EX.scala 30:24]
  wire [15:0] alu_io_restoration_pc; // @[EX.scala 30:24]
  wire [15:0] alu_io_rd_out; // @[EX.scala 30:24]
  wire [15:0] alu_io_pc_out; // @[EX.scala 30:24]
  wire  alu_io_mispredicted; // @[EX.scala 30:24]
  ALU alu ( // @[EX.scala 30:24]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_inst_info_valid(alu_io_inst_info_valid),
    .io_inst_info_rd_addr(alu_io_inst_info_rd_addr),
    .io_inst_info_rob_addr(alu_io_inst_info_rob_addr),
    .io_inst_info_ctrl_alu_op(alu_io_inst_info_ctrl_alu_op),
    .io_inst_info_ctrl_is_branch(alu_io_inst_info_ctrl_is_branch),
    .io_inst_info_ctrl_rf_w(alu_io_inst_info_ctrl_rf_w),
    .io_inst_info_ctrl_mem_r(alu_io_inst_info_ctrl_mem_r),
    .io_inst_info_ctrl_mem_w(alu_io_inst_info_ctrl_mem_w),
    .io_source_0(alu_io_source_0),
    .io_source_1(alu_io_source_1),
    .io_next_pc(alu_io_next_pc),
    .io_branch_pc(alu_io_branch_pc),
    .io_rd(alu_io_rd),
    .io_predict(alu_io_predict),
    .io_pc(alu_io_pc),
    .io_alu_out(alu_io_alu_out),
    .io_inst_info_out_valid(alu_io_inst_info_out_valid),
    .io_inst_info_out_rd_addr(alu_io_inst_info_out_rd_addr),
    .io_inst_info_out_rob_addr(alu_io_inst_info_out_rob_addr),
    .io_inst_info_out_ctrl_is_branch(alu_io_inst_info_out_ctrl_is_branch),
    .io_inst_info_out_ctrl_rf_w(alu_io_inst_info_out_ctrl_rf_w),
    .io_inst_info_out_ctrl_mem_r(alu_io_inst_info_out_ctrl_mem_r),
    .io_inst_info_out_ctrl_mem_w(alu_io_inst_info_out_ctrl_mem_w),
    .io_restoration_pc(alu_io_restoration_pc),
    .io_rd_out(alu_io_rd_out),
    .io_pc_out(alu_io_pc_out),
    .io_mispredicted(alu_io_mispredicted)
  );
  assign io_alu_out = alu_io_alu_out; // @[EX.scala 40:14]
  assign io_inst_info_out_valid = alu_io_inst_info_out_valid; // @[EX.scala 41:20]
  assign io_inst_info_out_rd_addr = alu_io_inst_info_out_rd_addr; // @[EX.scala 41:20]
  assign io_inst_info_out_rob_addr = alu_io_inst_info_out_rob_addr; // @[EX.scala 41:20]
  assign io_inst_info_out_ctrl_is_branch = alu_io_inst_info_out_ctrl_is_branch; // @[EX.scala 41:20]
  assign io_inst_info_out_ctrl_rf_w = alu_io_inst_info_out_ctrl_rf_w; // @[EX.scala 41:20]
  assign io_inst_info_out_ctrl_mem_r = alu_io_inst_info_out_ctrl_mem_r; // @[EX.scala 41:20]
  assign io_inst_info_out_ctrl_mem_w = alu_io_inst_info_out_ctrl_mem_w; // @[EX.scala 41:20]
  assign io_restoration_pc_out = alu_io_restoration_pc; // @[EX.scala 42:25]
  assign io_rd_out = alu_io_rd_out; // @[EX.scala 43:13]
  assign io_pc_out = alu_io_pc_out; // @[EX.scala 44:13]
  assign io_mispredicted = alu_io_mispredicted; // @[EX.scala 45:19]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_inst_info_valid = io_inst_info_valid; // @[EX.scala 31:20]
  assign alu_io_inst_info_rd_addr = io_inst_info_rd_addr; // @[EX.scala 31:20]
  assign alu_io_inst_info_rob_addr = io_inst_info_rob_addr; // @[EX.scala 31:20]
  assign alu_io_inst_info_ctrl_alu_op = io_inst_info_ctrl_alu_op; // @[EX.scala 31:20]
  assign alu_io_inst_info_ctrl_is_branch = io_inst_info_ctrl_is_branch; // @[EX.scala 31:20]
  assign alu_io_inst_info_ctrl_rf_w = io_inst_info_ctrl_rf_w; // @[EX.scala 31:20]
  assign alu_io_inst_info_ctrl_mem_r = io_inst_info_ctrl_mem_r; // @[EX.scala 31:20]
  assign alu_io_inst_info_ctrl_mem_w = io_inst_info_ctrl_mem_w; // @[EX.scala 31:20]
  assign alu_io_source_0 = io_source_0; // @[EX.scala 32:17]
  assign alu_io_source_1 = io_source_1; // @[EX.scala 32:17]
  assign alu_io_next_pc = io_next_pc; // @[EX.scala 33:18]
  assign alu_io_branch_pc = io_branch_pc; // @[EX.scala 34:20]
  assign alu_io_rd = io_rd; // @[EX.scala 35:13]
  assign alu_io_predict = io_predict; // @[EX.scala 36:18]
  assign alu_io_pc = io_pc; // @[EX.scala 37:13]
endmodule
module IM(
  input         clock,
  input         io_inst_info_valid,
  input  [2:0]  io_inst_info_rd_addr,
  input  [3:0]  io_inst_info_rob_addr,
  input         io_inst_info_ctrl_rf_w,
  input         io_inst_info_ctrl_mem_r,
  input         io_inst_info_ctrl_mem_w,
  input  [3:0]  io_rd_out,
  input  [3:0]  io_alu_out,
  output [15:0] io_mem_out
);
  reg [15:0] mem [0:127]; // @[IM.scala 18:27]
  reg [31:0] _RAND_0;
  wire [15:0] mem__T_1_data; // @[IM.scala 18:27]
  wire [6:0] mem__T_1_addr; // @[IM.scala 18:27]
  wire [15:0] mem__T_data; // @[IM.scala 18:27]
  wire [6:0] mem__T_addr; // @[IM.scala 18:27]
  wire  mem__T_mask; // @[IM.scala 18:27]
  wire  mem__T_en; // @[IM.scala 18:27]
  reg [15:0] out_data; // @[IM.scala 19:27]
  reg [31:0] _RAND_1;
  assign mem__T_1_addr = {{3'd0}, io_alu_out};
  assign mem__T_1_data = mem[mem__T_1_addr]; // @[IM.scala 18:27]
  assign mem__T_data = {{12'd0}, io_rd_out};
  assign mem__T_addr = {{3'd0}, io_alu_out};
  assign mem__T_mask = 1'h1;
  assign mem__T_en = io_inst_info_ctrl_mem_w;
  assign io_mem_out = out_data; // @[IM.scala 28:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_data = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_en & mem__T_mask) begin
      mem[mem__T_addr] <= mem__T_data; // @[IM.scala 18:27]
    end
    if (io_inst_info_ctrl_mem_w) begin
      out_data <= 16'h0;
    end else if (io_inst_info_ctrl_mem_r) begin
      out_data <= mem__T_1_data;
    end else begin
      out_data <= 16'h0;
    end
  end
endmodule
module ROB(
  input         clock,
  input         reset,
  input         io_used_num,
  input         io_graduate_0_valid,
  input  [15:0] io_graduate_0_bits_data,
  input  [2:0]  io_graduate_0_bits_inst_info_rd_addr,
  input         io_graduate_0_bits_inst_info_ctrl_rf_w,
  input  [3:0]  io_graduate_0_bits_addr,
  input         io_graduate_0_bits_mispredicted,
  input         io_graduate_1_valid,
  input  [15:0] io_graduate_1_bits_data,
  input  [2:0]  io_graduate_1_bits_inst_info_rd_addr,
  input         io_graduate_1_bits_inst_info_ctrl_rf_w,
  input  [3:0]  io_graduate_1_bits_addr,
  output [2:0]  io_commit_0_rd_addr,
  output        io_commit_0_rf_w,
  output [15:0] io_commit_0_data,
  output        io_unreserved_head_0_valid,
  output [3:0]  io_unreserved_head_0_bits
);
  reg [15:0] buf_0_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_0;
  reg [2:0] buf_0_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_1;
  reg  buf_0_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_2;
  reg  buf_0_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_3;
  reg  buf_0_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_4;
  reg [15:0] buf_1_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_5;
  reg [2:0] buf_1_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_6;
  reg  buf_1_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_7;
  reg  buf_1_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_8;
  reg  buf_1_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_9;
  reg [15:0] buf_2_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_10;
  reg [2:0] buf_2_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_11;
  reg  buf_2_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_12;
  reg  buf_2_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_13;
  reg  buf_2_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_14;
  reg [15:0] buf_3_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_15;
  reg [2:0] buf_3_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_16;
  reg  buf_3_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_17;
  reg  buf_3_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_18;
  reg  buf_3_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_19;
  reg [15:0] buf_4_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_20;
  reg [2:0] buf_4_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_21;
  reg  buf_4_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_22;
  reg  buf_4_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_23;
  reg  buf_4_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_24;
  reg [15:0] buf_5_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_25;
  reg [2:0] buf_5_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_26;
  reg  buf_5_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_27;
  reg  buf_5_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_28;
  reg  buf_5_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_29;
  reg [15:0] buf_6_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_30;
  reg [2:0] buf_6_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_31;
  reg  buf_6_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_32;
  reg  buf_6_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_33;
  reg  buf_6_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_34;
  reg [15:0] buf_7_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_35;
  reg [2:0] buf_7_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_36;
  reg  buf_7_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_37;
  reg  buf_7_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_38;
  reg  buf_7_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_39;
  reg [15:0] buf_8_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_40;
  reg [2:0] buf_8_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_41;
  reg  buf_8_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_42;
  reg  buf_8_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_43;
  reg  buf_8_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_44;
  reg [15:0] buf_9_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_45;
  reg [2:0] buf_9_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_46;
  reg  buf_9_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_47;
  reg  buf_9_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_48;
  reg  buf_9_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_49;
  reg [15:0] buf_10_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_50;
  reg [2:0] buf_10_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_51;
  reg  buf_10_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_52;
  reg  buf_10_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_53;
  reg  buf_10_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_54;
  reg [15:0] buf_11_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_55;
  reg [2:0] buf_11_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_56;
  reg  buf_11_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_57;
  reg  buf_11_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_58;
  reg  buf_11_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_59;
  reg [15:0] buf_12_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_60;
  reg [2:0] buf_12_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_61;
  reg  buf_12_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_62;
  reg  buf_12_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_63;
  reg  buf_12_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_64;
  reg [15:0] buf_13_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_65;
  reg [2:0] buf_13_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_66;
  reg  buf_13_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_67;
  reg  buf_13_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_68;
  reg  buf_13_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_69;
  reg [15:0] buf_14_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_70;
  reg [2:0] buf_14_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_71;
  reg  buf_14_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_72;
  reg  buf_14_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_73;
  reg  buf_14_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_74;
  reg [15:0] buf_15_data; // @[ROB.scala 40:35]
  reg [31:0] _RAND_75;
  reg [2:0] buf_15_inst_info_rd_addr; // @[ROB.scala 40:35]
  reg [31:0] _RAND_76;
  reg  buf_15_inst_info_ctrl_rf_w; // @[ROB.scala 40:35]
  reg [31:0] _RAND_77;
  reg  buf_15_reserved; // @[ROB.scala 40:35]
  reg [31:0] _RAND_78;
  reg  buf_15_committable; // @[ROB.scala 40:35]
  reg [31:0] _RAND_79;
  reg [3:0] uncommited; // @[ROB.scala 42:33]
  reg [31:0] _RAND_80;
  wire [4:0] _T_3; // @[ROB.scala 44:48]
  wire [3:0] _T_4; // @[ROB.scala 44:48]
  wire [15:0] _GEN_16; // @[ROB.scala 43:50]
  wire [2:0] _GEN_20; // @[ROB.scala 43:50]
  wire  _GEN_25; // @[ROB.scala 43:50]
  wire  _GEN_31; // @[ROB.scala 43:50]
  wire [15:0] _GEN_32; // @[ROB.scala 43:50]
  wire [2:0] _GEN_36; // @[ROB.scala 43:50]
  wire  _GEN_41; // @[ROB.scala 43:50]
  wire  _GEN_47; // @[ROB.scala 43:50]
  wire [15:0] _GEN_48; // @[ROB.scala 43:50]
  wire [2:0] _GEN_52; // @[ROB.scala 43:50]
  wire  _GEN_57; // @[ROB.scala 43:50]
  wire  _GEN_63; // @[ROB.scala 43:50]
  wire [15:0] _GEN_64; // @[ROB.scala 43:50]
  wire [2:0] _GEN_68; // @[ROB.scala 43:50]
  wire  _GEN_73; // @[ROB.scala 43:50]
  wire  _GEN_79; // @[ROB.scala 43:50]
  wire [15:0] _GEN_80; // @[ROB.scala 43:50]
  wire [2:0] _GEN_84; // @[ROB.scala 43:50]
  wire  _GEN_89; // @[ROB.scala 43:50]
  wire  _GEN_95; // @[ROB.scala 43:50]
  wire [15:0] _GEN_96; // @[ROB.scala 43:50]
  wire [2:0] _GEN_100; // @[ROB.scala 43:50]
  wire  _GEN_105; // @[ROB.scala 43:50]
  wire  _GEN_111; // @[ROB.scala 43:50]
  wire [15:0] _GEN_112; // @[ROB.scala 43:50]
  wire [2:0] _GEN_116; // @[ROB.scala 43:50]
  wire  _GEN_121; // @[ROB.scala 43:50]
  wire  _GEN_127; // @[ROB.scala 43:50]
  wire [15:0] _GEN_128; // @[ROB.scala 43:50]
  wire [2:0] _GEN_132; // @[ROB.scala 43:50]
  wire  _GEN_137; // @[ROB.scala 43:50]
  wire  _GEN_143; // @[ROB.scala 43:50]
  wire [15:0] _GEN_144; // @[ROB.scala 43:50]
  wire [2:0] _GEN_148; // @[ROB.scala 43:50]
  wire  _GEN_153; // @[ROB.scala 43:50]
  wire  _GEN_159; // @[ROB.scala 43:50]
  wire [15:0] _GEN_160; // @[ROB.scala 43:50]
  wire [2:0] _GEN_164; // @[ROB.scala 43:50]
  wire  _GEN_169; // @[ROB.scala 43:50]
  wire  _GEN_175; // @[ROB.scala 43:50]
  wire [15:0] _GEN_176; // @[ROB.scala 43:50]
  wire [2:0] _GEN_180; // @[ROB.scala 43:50]
  wire  _GEN_185; // @[ROB.scala 43:50]
  wire  _GEN_191; // @[ROB.scala 43:50]
  wire [15:0] _GEN_192; // @[ROB.scala 43:50]
  wire [2:0] _GEN_196; // @[ROB.scala 43:50]
  wire  _GEN_201; // @[ROB.scala 43:50]
  wire  _GEN_207; // @[ROB.scala 43:50]
  wire [15:0] _GEN_208; // @[ROB.scala 43:50]
  wire [2:0] _GEN_212; // @[ROB.scala 43:50]
  wire  _GEN_217; // @[ROB.scala 43:50]
  wire  _GEN_223; // @[ROB.scala 43:50]
  wire [15:0] _GEN_224; // @[ROB.scala 43:50]
  wire [2:0] _GEN_228; // @[ROB.scala 43:50]
  wire  _GEN_233; // @[ROB.scala 43:50]
  wire  _GEN_239; // @[ROB.scala 43:50]
  wire [15:0] _GEN_240; // @[ROB.scala 43:50]
  wire [2:0] _GEN_244; // @[ROB.scala 43:50]
  wire  _GEN_249; // @[ROB.scala 43:50]
  wire  commitable_0; // @[ROB.scala 43:50]
  wire [3:0] _GEN_1571; // @[ROB.scala 50:41]
  wire [3:0] next_uncommited; // @[ROB.scala 50:41]
  wire  _T_7; // @[ROB.scala 53:136]
  wire  _T_8_valid; // @[ROB.scala 53:126]
  wire [3:0] _T_8_bits_addr; // @[ROB.scala 53:126]
  wire  _T_8_bits_mispredicted; // @[ROB.scala 53:126]
  wire  mispredicted; // @[ROB.scala 54:53]
  reg [3:0] unreserved; // @[ROB.scala 57:33]
  reg [31:0] _RAND_81;
  wire [3:0] _GEN_1572; // @[ROB.scala 58:46]
  wire [3:0] unreserved_add_used; // @[ROB.scala 58:46]
  wire  _GEN_286; // @[ROB.scala 59:41]
  wire  _GEN_302; // @[ROB.scala 59:41]
  wire  _GEN_318; // @[ROB.scala 59:41]
  wire  _GEN_334; // @[ROB.scala 59:41]
  wire  _GEN_350; // @[ROB.scala 59:41]
  wire  _GEN_366; // @[ROB.scala 59:41]
  wire  _GEN_382; // @[ROB.scala 59:41]
  wire  _GEN_398; // @[ROB.scala 59:41]
  wire  _GEN_414; // @[ROB.scala 59:41]
  wire  _GEN_430; // @[ROB.scala 59:41]
  wire  _GEN_446; // @[ROB.scala 59:41]
  wire  _GEN_462; // @[ROB.scala 59:41]
  wire  _GEN_478; // @[ROB.scala 59:41]
  wire  _GEN_494; // @[ROB.scala 59:41]
  wire  _GEN_510; // @[ROB.scala 59:41]
  wire  unreserved_add_used_valid; // @[ROB.scala 59:41]
  wire [3:0] _T_11; // @[Mux.scala 87:16]
  wire [3:0] next_unreserved; // @[Mux.scala 87:16]
  wire  _T_12; // @[ROB.scala 68:36]
  wire  _T_13; // @[ROB.scala 68:20]
  wire  _T_14_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_14_bits_addr; // @[ROB.scala 68:10]
  wire  _T_16; // @[ROB.scala 71:27]
  wire  _T_17; // @[ROB.scala 71:61]
  wire  _T_18; // @[ROB.scala 71:41]
  wire  _T_19; // @[ROB.scala 71:75]
  wire  _T_20; // @[ROB.scala 71:68]
  wire  _T_21; // @[ROB.scala 72:27]
  wire  _T_24; // @[ROB.scala 72:61]
  wire  _T_25; // @[ROB.scala 72:40]
  wire  _T_26; // @[ROB.scala 71:89]
  wire  _T_27; // @[ROB.scala 70:56]
  wire  _T_28; // @[ROB.scala 74:25]
  wire  _T_29; // @[ROB.scala 75:20]
  wire  _T_30; // @[ROB.scala 75:55]
  wire  _T_31; // @[ROB.scala 75:69]
  wire  _T_32; // @[ROB.scala 75:62]
  wire  _T_33; // @[ROB.scala 75:40]
  wire  _T_34; // @[ROB.scala 76:20]
  wire  _T_37; // @[ROB.scala 76:65]
  wire  _T_38; // @[ROB.scala 76:39]
  wire  _T_39; // @[ROB.scala 75:89]
  wire  _T_40; // @[ROB.scala 74:39]
  wire  _T_41; // @[ROB.scala 79:20]
  wire  _T_42; // @[ROB.scala 79:55]
  wire  _T_43; // @[ROB.scala 79:69]
  wire  _T_44; // @[ROB.scala 79:62]
  wire  _T_45; // @[ROB.scala 79:40]
  wire  _T_46; // @[ROB.scala 80:20]
  wire  _T_49; // @[ROB.scala 80:66]
  wire  _T_50; // @[ROB.scala 80:40]
  wire  _T_51; // @[ROB.scala 79:89]
  wire  _T_52; // @[ROB.scala 82:60]
  wire  _T_53; // @[ROB.scala 82:38]
  wire  _GEN_512; // @[ROB.scala 98:31]
  wire  _GEN_513; // @[ROB.scala 98:31]
  wire  _GEN_514; // @[ROB.scala 94:29]
  wire  _GEN_529; // @[ROB.scala 94:29]
  wire  _GEN_530; // @[ROB.scala 92:32]
  wire  _T_54; // @[ROB.scala 68:36]
  wire  _T_55; // @[ROB.scala 68:20]
  wire  _T_56_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_56_bits_addr; // @[ROB.scala 68:10]
  wire  _T_59; // @[ROB.scala 71:61]
  wire  _T_60; // @[ROB.scala 71:41]
  wire  _T_61; // @[ROB.scala 71:75]
  wire  _T_62; // @[ROB.scala 71:68]
  wire  _T_66; // @[ROB.scala 72:61]
  wire  _T_67; // @[ROB.scala 72:40]
  wire  _T_68; // @[ROB.scala 71:89]
  wire  _T_69; // @[ROB.scala 70:56]
  wire  _T_72; // @[ROB.scala 75:55]
  wire  _T_73; // @[ROB.scala 75:69]
  wire  _T_74; // @[ROB.scala 75:62]
  wire  _T_75; // @[ROB.scala 75:40]
  wire  _T_79; // @[ROB.scala 76:65]
  wire  _T_80; // @[ROB.scala 76:39]
  wire  _T_81; // @[ROB.scala 75:89]
  wire  _T_82; // @[ROB.scala 74:39]
  wire  _T_84; // @[ROB.scala 79:55]
  wire  _T_85; // @[ROB.scala 79:69]
  wire  _T_86; // @[ROB.scala 79:62]
  wire  _T_87; // @[ROB.scala 79:40]
  wire  _T_91; // @[ROB.scala 80:66]
  wire  _T_92; // @[ROB.scala 80:40]
  wire  _T_93; // @[ROB.scala 79:89]
  wire  _T_94; // @[ROB.scala 82:60]
  wire  _T_95; // @[ROB.scala 82:38]
  wire  _GEN_562; // @[ROB.scala 98:31]
  wire  _GEN_563; // @[ROB.scala 98:31]
  wire  _GEN_564; // @[ROB.scala 94:29]
  wire  _GEN_579; // @[ROB.scala 94:29]
  wire  _GEN_580; // @[ROB.scala 92:32]
  wire  _T_96; // @[ROB.scala 68:36]
  wire  _T_97; // @[ROB.scala 68:20]
  wire  _T_98_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_98_bits_addr; // @[ROB.scala 68:10]
  wire  _T_101; // @[ROB.scala 71:61]
  wire  _T_102; // @[ROB.scala 71:41]
  wire  _T_103; // @[ROB.scala 71:75]
  wire  _T_104; // @[ROB.scala 71:68]
  wire  _T_108; // @[ROB.scala 72:61]
  wire  _T_109; // @[ROB.scala 72:40]
  wire  _T_110; // @[ROB.scala 71:89]
  wire  _T_111; // @[ROB.scala 70:56]
  wire  _T_114; // @[ROB.scala 75:55]
  wire  _T_115; // @[ROB.scala 75:69]
  wire  _T_116; // @[ROB.scala 75:62]
  wire  _T_117; // @[ROB.scala 75:40]
  wire  _T_121; // @[ROB.scala 76:65]
  wire  _T_122; // @[ROB.scala 76:39]
  wire  _T_123; // @[ROB.scala 75:89]
  wire  _T_124; // @[ROB.scala 74:39]
  wire  _T_126; // @[ROB.scala 79:55]
  wire  _T_127; // @[ROB.scala 79:69]
  wire  _T_128; // @[ROB.scala 79:62]
  wire  _T_129; // @[ROB.scala 79:40]
  wire  _T_133; // @[ROB.scala 80:66]
  wire  _T_134; // @[ROB.scala 80:40]
  wire  _T_135; // @[ROB.scala 79:89]
  wire  _T_136; // @[ROB.scala 82:60]
  wire  _T_137; // @[ROB.scala 82:38]
  wire  _GEN_612; // @[ROB.scala 98:31]
  wire  _GEN_613; // @[ROB.scala 98:31]
  wire  _GEN_614; // @[ROB.scala 94:29]
  wire  _GEN_629; // @[ROB.scala 94:29]
  wire  _GEN_630; // @[ROB.scala 92:32]
  wire  _T_138; // @[ROB.scala 68:36]
  wire  _T_139; // @[ROB.scala 68:20]
  wire  _T_140_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_140_bits_addr; // @[ROB.scala 68:10]
  wire  _T_143; // @[ROB.scala 71:61]
  wire  _T_144; // @[ROB.scala 71:41]
  wire  _T_145; // @[ROB.scala 71:75]
  wire  _T_146; // @[ROB.scala 71:68]
  wire  _T_150; // @[ROB.scala 72:61]
  wire  _T_151; // @[ROB.scala 72:40]
  wire  _T_152; // @[ROB.scala 71:89]
  wire  _T_153; // @[ROB.scala 70:56]
  wire  _T_156; // @[ROB.scala 75:55]
  wire  _T_157; // @[ROB.scala 75:69]
  wire  _T_158; // @[ROB.scala 75:62]
  wire  _T_159; // @[ROB.scala 75:40]
  wire  _T_163; // @[ROB.scala 76:65]
  wire  _T_164; // @[ROB.scala 76:39]
  wire  _T_165; // @[ROB.scala 75:89]
  wire  _T_166; // @[ROB.scala 74:39]
  wire  _T_168; // @[ROB.scala 79:55]
  wire  _T_169; // @[ROB.scala 79:69]
  wire  _T_170; // @[ROB.scala 79:62]
  wire  _T_171; // @[ROB.scala 79:40]
  wire  _T_175; // @[ROB.scala 80:66]
  wire  _T_176; // @[ROB.scala 80:40]
  wire  _T_177; // @[ROB.scala 79:89]
  wire  _T_178; // @[ROB.scala 82:60]
  wire  _T_179; // @[ROB.scala 82:38]
  wire  _GEN_662; // @[ROB.scala 98:31]
  wire  _GEN_663; // @[ROB.scala 98:31]
  wire  _GEN_664; // @[ROB.scala 94:29]
  wire  _GEN_679; // @[ROB.scala 94:29]
  wire  _GEN_680; // @[ROB.scala 92:32]
  wire  _T_180; // @[ROB.scala 68:36]
  wire  _T_181; // @[ROB.scala 68:20]
  wire  _T_182_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_182_bits_addr; // @[ROB.scala 68:10]
  wire  _T_185; // @[ROB.scala 71:61]
  wire  _T_186; // @[ROB.scala 71:41]
  wire  _T_187; // @[ROB.scala 71:75]
  wire  _T_188; // @[ROB.scala 71:68]
  wire  _T_192; // @[ROB.scala 72:61]
  wire  _T_193; // @[ROB.scala 72:40]
  wire  _T_194; // @[ROB.scala 71:89]
  wire  _T_195; // @[ROB.scala 70:56]
  wire  _T_198; // @[ROB.scala 75:55]
  wire  _T_199; // @[ROB.scala 75:69]
  wire  _T_200; // @[ROB.scala 75:62]
  wire  _T_201; // @[ROB.scala 75:40]
  wire  _T_205; // @[ROB.scala 76:65]
  wire  _T_206; // @[ROB.scala 76:39]
  wire  _T_207; // @[ROB.scala 75:89]
  wire  _T_208; // @[ROB.scala 74:39]
  wire  _T_210; // @[ROB.scala 79:55]
  wire  _T_211; // @[ROB.scala 79:69]
  wire  _T_212; // @[ROB.scala 79:62]
  wire  _T_213; // @[ROB.scala 79:40]
  wire  _T_217; // @[ROB.scala 80:66]
  wire  _T_218; // @[ROB.scala 80:40]
  wire  _T_219; // @[ROB.scala 79:89]
  wire  _T_220; // @[ROB.scala 82:60]
  wire  _T_221; // @[ROB.scala 82:38]
  wire  _GEN_712; // @[ROB.scala 98:31]
  wire  _GEN_713; // @[ROB.scala 98:31]
  wire  _GEN_714; // @[ROB.scala 94:29]
  wire  _GEN_729; // @[ROB.scala 94:29]
  wire  _GEN_730; // @[ROB.scala 92:32]
  wire  _T_222; // @[ROB.scala 68:36]
  wire  _T_223; // @[ROB.scala 68:20]
  wire  _T_224_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_224_bits_addr; // @[ROB.scala 68:10]
  wire  _T_227; // @[ROB.scala 71:61]
  wire  _T_228; // @[ROB.scala 71:41]
  wire  _T_229; // @[ROB.scala 71:75]
  wire  _T_230; // @[ROB.scala 71:68]
  wire  _T_234; // @[ROB.scala 72:61]
  wire  _T_235; // @[ROB.scala 72:40]
  wire  _T_236; // @[ROB.scala 71:89]
  wire  _T_237; // @[ROB.scala 70:56]
  wire  _T_240; // @[ROB.scala 75:55]
  wire  _T_241; // @[ROB.scala 75:69]
  wire  _T_242; // @[ROB.scala 75:62]
  wire  _T_243; // @[ROB.scala 75:40]
  wire  _T_247; // @[ROB.scala 76:65]
  wire  _T_248; // @[ROB.scala 76:39]
  wire  _T_249; // @[ROB.scala 75:89]
  wire  _T_250; // @[ROB.scala 74:39]
  wire  _T_252; // @[ROB.scala 79:55]
  wire  _T_253; // @[ROB.scala 79:69]
  wire  _T_254; // @[ROB.scala 79:62]
  wire  _T_255; // @[ROB.scala 79:40]
  wire  _T_259; // @[ROB.scala 80:66]
  wire  _T_260; // @[ROB.scala 80:40]
  wire  _T_261; // @[ROB.scala 79:89]
  wire  _T_262; // @[ROB.scala 82:60]
  wire  _T_263; // @[ROB.scala 82:38]
  wire  _GEN_762; // @[ROB.scala 98:31]
  wire  _GEN_763; // @[ROB.scala 98:31]
  wire  _GEN_764; // @[ROB.scala 94:29]
  wire  _GEN_779; // @[ROB.scala 94:29]
  wire  _GEN_780; // @[ROB.scala 92:32]
  wire  _T_264; // @[ROB.scala 68:36]
  wire  _T_265; // @[ROB.scala 68:20]
  wire  _T_266_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_266_bits_addr; // @[ROB.scala 68:10]
  wire  _T_269; // @[ROB.scala 71:61]
  wire  _T_270; // @[ROB.scala 71:41]
  wire  _T_271; // @[ROB.scala 71:75]
  wire  _T_272; // @[ROB.scala 71:68]
  wire  _T_276; // @[ROB.scala 72:61]
  wire  _T_277; // @[ROB.scala 72:40]
  wire  _T_278; // @[ROB.scala 71:89]
  wire  _T_279; // @[ROB.scala 70:56]
  wire  _T_282; // @[ROB.scala 75:55]
  wire  _T_283; // @[ROB.scala 75:69]
  wire  _T_284; // @[ROB.scala 75:62]
  wire  _T_285; // @[ROB.scala 75:40]
  wire  _T_289; // @[ROB.scala 76:65]
  wire  _T_290; // @[ROB.scala 76:39]
  wire  _T_291; // @[ROB.scala 75:89]
  wire  _T_292; // @[ROB.scala 74:39]
  wire  _T_294; // @[ROB.scala 79:55]
  wire  _T_295; // @[ROB.scala 79:69]
  wire  _T_296; // @[ROB.scala 79:62]
  wire  _T_297; // @[ROB.scala 79:40]
  wire  _T_301; // @[ROB.scala 80:66]
  wire  _T_302; // @[ROB.scala 80:40]
  wire  _T_303; // @[ROB.scala 79:89]
  wire  _T_304; // @[ROB.scala 82:60]
  wire  _T_305; // @[ROB.scala 82:38]
  wire  _GEN_812; // @[ROB.scala 98:31]
  wire  _GEN_813; // @[ROB.scala 98:31]
  wire  _GEN_814; // @[ROB.scala 94:29]
  wire  _GEN_829; // @[ROB.scala 94:29]
  wire  _GEN_830; // @[ROB.scala 92:32]
  wire  _T_306; // @[ROB.scala 68:36]
  wire  _T_307; // @[ROB.scala 68:20]
  wire  _T_308_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_308_bits_addr; // @[ROB.scala 68:10]
  wire  _T_311; // @[ROB.scala 71:61]
  wire  _T_312; // @[ROB.scala 71:41]
  wire  _T_313; // @[ROB.scala 71:75]
  wire  _T_314; // @[ROB.scala 71:68]
  wire  _T_318; // @[ROB.scala 72:61]
  wire  _T_319; // @[ROB.scala 72:40]
  wire  _T_320; // @[ROB.scala 71:89]
  wire  _T_321; // @[ROB.scala 70:56]
  wire  _T_324; // @[ROB.scala 75:55]
  wire  _T_325; // @[ROB.scala 75:69]
  wire  _T_326; // @[ROB.scala 75:62]
  wire  _T_327; // @[ROB.scala 75:40]
  wire  _T_331; // @[ROB.scala 76:65]
  wire  _T_332; // @[ROB.scala 76:39]
  wire  _T_333; // @[ROB.scala 75:89]
  wire  _T_334; // @[ROB.scala 74:39]
  wire  _T_336; // @[ROB.scala 79:55]
  wire  _T_337; // @[ROB.scala 79:69]
  wire  _T_338; // @[ROB.scala 79:62]
  wire  _T_339; // @[ROB.scala 79:40]
  wire  _T_343; // @[ROB.scala 80:66]
  wire  _T_344; // @[ROB.scala 80:40]
  wire  _T_345; // @[ROB.scala 79:89]
  wire  _T_346; // @[ROB.scala 82:60]
  wire  _T_347; // @[ROB.scala 82:38]
  wire  _GEN_862; // @[ROB.scala 98:31]
  wire  _GEN_863; // @[ROB.scala 98:31]
  wire  _GEN_864; // @[ROB.scala 94:29]
  wire  _GEN_879; // @[ROB.scala 94:29]
  wire  _GEN_880; // @[ROB.scala 92:32]
  wire  _T_348; // @[ROB.scala 68:36]
  wire  _T_349; // @[ROB.scala 68:20]
  wire  _T_350_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_350_bits_addr; // @[ROB.scala 68:10]
  wire  _T_353; // @[ROB.scala 71:61]
  wire  _T_354; // @[ROB.scala 71:41]
  wire  _T_355; // @[ROB.scala 71:75]
  wire  _T_356; // @[ROB.scala 71:68]
  wire  _T_360; // @[ROB.scala 72:61]
  wire  _T_361; // @[ROB.scala 72:40]
  wire  _T_362; // @[ROB.scala 71:89]
  wire  _T_363; // @[ROB.scala 70:56]
  wire  _T_366; // @[ROB.scala 75:55]
  wire  _T_367; // @[ROB.scala 75:69]
  wire  _T_368; // @[ROB.scala 75:62]
  wire  _T_369; // @[ROB.scala 75:40]
  wire  _T_373; // @[ROB.scala 76:65]
  wire  _T_374; // @[ROB.scala 76:39]
  wire  _T_375; // @[ROB.scala 75:89]
  wire  _T_376; // @[ROB.scala 74:39]
  wire  _T_378; // @[ROB.scala 79:55]
  wire  _T_379; // @[ROB.scala 79:69]
  wire  _T_380; // @[ROB.scala 79:62]
  wire  _T_381; // @[ROB.scala 79:40]
  wire  _T_385; // @[ROB.scala 80:66]
  wire  _T_386; // @[ROB.scala 80:40]
  wire  _T_387; // @[ROB.scala 79:89]
  wire  _T_388; // @[ROB.scala 82:60]
  wire  _T_389; // @[ROB.scala 82:38]
  wire  _GEN_912; // @[ROB.scala 98:31]
  wire  _GEN_913; // @[ROB.scala 98:31]
  wire  _GEN_914; // @[ROB.scala 94:29]
  wire  _GEN_929; // @[ROB.scala 94:29]
  wire  _GEN_930; // @[ROB.scala 92:32]
  wire  _T_390; // @[ROB.scala 68:36]
  wire  _T_391; // @[ROB.scala 68:20]
  wire  _T_392_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_392_bits_addr; // @[ROB.scala 68:10]
  wire  _T_395; // @[ROB.scala 71:61]
  wire  _T_396; // @[ROB.scala 71:41]
  wire  _T_397; // @[ROB.scala 71:75]
  wire  _T_398; // @[ROB.scala 71:68]
  wire  _T_402; // @[ROB.scala 72:61]
  wire  _T_403; // @[ROB.scala 72:40]
  wire  _T_404; // @[ROB.scala 71:89]
  wire  _T_405; // @[ROB.scala 70:56]
  wire  _T_408; // @[ROB.scala 75:55]
  wire  _T_409; // @[ROB.scala 75:69]
  wire  _T_410; // @[ROB.scala 75:62]
  wire  _T_411; // @[ROB.scala 75:40]
  wire  _T_415; // @[ROB.scala 76:65]
  wire  _T_416; // @[ROB.scala 76:39]
  wire  _T_417; // @[ROB.scala 75:89]
  wire  _T_418; // @[ROB.scala 74:39]
  wire  _T_420; // @[ROB.scala 79:55]
  wire  _T_421; // @[ROB.scala 79:69]
  wire  _T_422; // @[ROB.scala 79:62]
  wire  _T_423; // @[ROB.scala 79:40]
  wire  _T_427; // @[ROB.scala 80:66]
  wire  _T_428; // @[ROB.scala 80:40]
  wire  _T_429; // @[ROB.scala 79:89]
  wire  _T_430; // @[ROB.scala 82:60]
  wire  _T_431; // @[ROB.scala 82:38]
  wire  _GEN_962; // @[ROB.scala 98:31]
  wire  _GEN_963; // @[ROB.scala 98:31]
  wire  _GEN_964; // @[ROB.scala 94:29]
  wire  _GEN_979; // @[ROB.scala 94:29]
  wire  _GEN_980; // @[ROB.scala 92:32]
  wire  _T_432; // @[ROB.scala 68:36]
  wire  _T_433; // @[ROB.scala 68:20]
  wire  _T_434_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_434_bits_addr; // @[ROB.scala 68:10]
  wire  _T_437; // @[ROB.scala 71:61]
  wire  _T_438; // @[ROB.scala 71:41]
  wire  _T_439; // @[ROB.scala 71:75]
  wire  _T_440; // @[ROB.scala 71:68]
  wire  _T_444; // @[ROB.scala 72:61]
  wire  _T_445; // @[ROB.scala 72:40]
  wire  _T_446; // @[ROB.scala 71:89]
  wire  _T_447; // @[ROB.scala 70:56]
  wire  _T_450; // @[ROB.scala 75:55]
  wire  _T_451; // @[ROB.scala 75:69]
  wire  _T_452; // @[ROB.scala 75:62]
  wire  _T_453; // @[ROB.scala 75:40]
  wire  _T_457; // @[ROB.scala 76:65]
  wire  _T_458; // @[ROB.scala 76:39]
  wire  _T_459; // @[ROB.scala 75:89]
  wire  _T_460; // @[ROB.scala 74:39]
  wire  _T_462; // @[ROB.scala 79:55]
  wire  _T_463; // @[ROB.scala 79:69]
  wire  _T_464; // @[ROB.scala 79:62]
  wire  _T_465; // @[ROB.scala 79:40]
  wire  _T_469; // @[ROB.scala 80:66]
  wire  _T_470; // @[ROB.scala 80:40]
  wire  _T_471; // @[ROB.scala 79:89]
  wire  _T_472; // @[ROB.scala 82:60]
  wire  _T_473; // @[ROB.scala 82:38]
  wire  _GEN_1012; // @[ROB.scala 98:31]
  wire  _GEN_1013; // @[ROB.scala 98:31]
  wire  _GEN_1014; // @[ROB.scala 94:29]
  wire  _GEN_1029; // @[ROB.scala 94:29]
  wire  _GEN_1030; // @[ROB.scala 92:32]
  wire  _T_474; // @[ROB.scala 68:36]
  wire  _T_475; // @[ROB.scala 68:20]
  wire  _T_476_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_476_bits_addr; // @[ROB.scala 68:10]
  wire  _T_479; // @[ROB.scala 71:61]
  wire  _T_480; // @[ROB.scala 71:41]
  wire  _T_481; // @[ROB.scala 71:75]
  wire  _T_482; // @[ROB.scala 71:68]
  wire  _T_486; // @[ROB.scala 72:61]
  wire  _T_487; // @[ROB.scala 72:40]
  wire  _T_488; // @[ROB.scala 71:89]
  wire  _T_489; // @[ROB.scala 70:56]
  wire  _T_492; // @[ROB.scala 75:55]
  wire  _T_493; // @[ROB.scala 75:69]
  wire  _T_494; // @[ROB.scala 75:62]
  wire  _T_495; // @[ROB.scala 75:40]
  wire  _T_499; // @[ROB.scala 76:65]
  wire  _T_500; // @[ROB.scala 76:39]
  wire  _T_501; // @[ROB.scala 75:89]
  wire  _T_502; // @[ROB.scala 74:39]
  wire  _T_504; // @[ROB.scala 79:55]
  wire  _T_505; // @[ROB.scala 79:69]
  wire  _T_506; // @[ROB.scala 79:62]
  wire  _T_507; // @[ROB.scala 79:40]
  wire  _T_511; // @[ROB.scala 80:66]
  wire  _T_512; // @[ROB.scala 80:40]
  wire  _T_513; // @[ROB.scala 79:89]
  wire  _T_514; // @[ROB.scala 82:60]
  wire  _T_515; // @[ROB.scala 82:38]
  wire  _GEN_1062; // @[ROB.scala 98:31]
  wire  _GEN_1063; // @[ROB.scala 98:31]
  wire  _GEN_1064; // @[ROB.scala 94:29]
  wire  _GEN_1079; // @[ROB.scala 94:29]
  wire  _GEN_1080; // @[ROB.scala 92:32]
  wire  _T_516; // @[ROB.scala 68:36]
  wire  _T_517; // @[ROB.scala 68:20]
  wire  _T_518_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_518_bits_addr; // @[ROB.scala 68:10]
  wire  _T_521; // @[ROB.scala 71:61]
  wire  _T_522; // @[ROB.scala 71:41]
  wire  _T_523; // @[ROB.scala 71:75]
  wire  _T_524; // @[ROB.scala 71:68]
  wire  _T_528; // @[ROB.scala 72:61]
  wire  _T_529; // @[ROB.scala 72:40]
  wire  _T_530; // @[ROB.scala 71:89]
  wire  _T_531; // @[ROB.scala 70:56]
  wire  _T_534; // @[ROB.scala 75:55]
  wire  _T_535; // @[ROB.scala 75:69]
  wire  _T_536; // @[ROB.scala 75:62]
  wire  _T_537; // @[ROB.scala 75:40]
  wire  _T_541; // @[ROB.scala 76:65]
  wire  _T_542; // @[ROB.scala 76:39]
  wire  _T_543; // @[ROB.scala 75:89]
  wire  _T_544; // @[ROB.scala 74:39]
  wire  _T_546; // @[ROB.scala 79:55]
  wire  _T_547; // @[ROB.scala 79:69]
  wire  _T_548; // @[ROB.scala 79:62]
  wire  _T_549; // @[ROB.scala 79:40]
  wire  _T_553; // @[ROB.scala 80:66]
  wire  _T_554; // @[ROB.scala 80:40]
  wire  _T_555; // @[ROB.scala 79:89]
  wire  _T_556; // @[ROB.scala 82:60]
  wire  _T_557; // @[ROB.scala 82:38]
  wire  _GEN_1112; // @[ROB.scala 98:31]
  wire  _GEN_1113; // @[ROB.scala 98:31]
  wire  _GEN_1114; // @[ROB.scala 94:29]
  wire  _GEN_1129; // @[ROB.scala 94:29]
  wire  _GEN_1130; // @[ROB.scala 92:32]
  wire  _T_558; // @[ROB.scala 68:36]
  wire  _T_559; // @[ROB.scala 68:20]
  wire  _T_560_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_560_bits_addr; // @[ROB.scala 68:10]
  wire  _T_563; // @[ROB.scala 71:61]
  wire  _T_564; // @[ROB.scala 71:41]
  wire  _T_565; // @[ROB.scala 71:75]
  wire  _T_566; // @[ROB.scala 71:68]
  wire  _T_570; // @[ROB.scala 72:61]
  wire  _T_571; // @[ROB.scala 72:40]
  wire  _T_572; // @[ROB.scala 71:89]
  wire  _T_573; // @[ROB.scala 70:56]
  wire  _T_576; // @[ROB.scala 75:55]
  wire  _T_577; // @[ROB.scala 75:69]
  wire  _T_578; // @[ROB.scala 75:62]
  wire  _T_579; // @[ROB.scala 75:40]
  wire  _T_583; // @[ROB.scala 76:65]
  wire  _T_584; // @[ROB.scala 76:39]
  wire  _T_585; // @[ROB.scala 75:89]
  wire  _T_586; // @[ROB.scala 74:39]
  wire  _T_588; // @[ROB.scala 79:55]
  wire  _T_589; // @[ROB.scala 79:69]
  wire  _T_590; // @[ROB.scala 79:62]
  wire  _T_591; // @[ROB.scala 79:40]
  wire  _T_595; // @[ROB.scala 80:66]
  wire  _T_596; // @[ROB.scala 80:40]
  wire  _T_597; // @[ROB.scala 79:89]
  wire  _T_598; // @[ROB.scala 82:60]
  wire  _T_599; // @[ROB.scala 82:38]
  wire  _GEN_1162; // @[ROB.scala 98:31]
  wire  _GEN_1163; // @[ROB.scala 98:31]
  wire  _GEN_1164; // @[ROB.scala 94:29]
  wire  _GEN_1179; // @[ROB.scala 94:29]
  wire  _GEN_1180; // @[ROB.scala 92:32]
  wire  _T_600; // @[ROB.scala 68:36]
  wire  _T_601; // @[ROB.scala 68:20]
  wire  _T_602_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_602_bits_addr; // @[ROB.scala 68:10]
  wire  _T_605; // @[ROB.scala 71:61]
  wire  _T_606; // @[ROB.scala 71:41]
  wire  _T_607; // @[ROB.scala 71:75]
  wire  _T_608; // @[ROB.scala 71:68]
  wire  _T_612; // @[ROB.scala 72:61]
  wire  _T_613; // @[ROB.scala 72:40]
  wire  _T_614; // @[ROB.scala 71:89]
  wire  _T_615; // @[ROB.scala 70:56]
  wire  _T_618; // @[ROB.scala 75:55]
  wire  _T_619; // @[ROB.scala 75:69]
  wire  _T_620; // @[ROB.scala 75:62]
  wire  _T_621; // @[ROB.scala 75:40]
  wire  _T_625; // @[ROB.scala 76:65]
  wire  _T_626; // @[ROB.scala 76:39]
  wire  _T_627; // @[ROB.scala 75:89]
  wire  _T_628; // @[ROB.scala 74:39]
  wire  _T_630; // @[ROB.scala 79:55]
  wire  _T_631; // @[ROB.scala 79:69]
  wire  _T_632; // @[ROB.scala 79:62]
  wire  _T_633; // @[ROB.scala 79:40]
  wire  _T_637; // @[ROB.scala 80:66]
  wire  _T_638; // @[ROB.scala 80:40]
  wire  _T_639; // @[ROB.scala 79:89]
  wire  _T_640; // @[ROB.scala 82:60]
  wire  _T_641; // @[ROB.scala 82:38]
  wire  _GEN_1212; // @[ROB.scala 98:31]
  wire  _GEN_1213; // @[ROB.scala 98:31]
  wire  _GEN_1214; // @[ROB.scala 94:29]
  wire  _GEN_1229; // @[ROB.scala 94:29]
  wire  _GEN_1230; // @[ROB.scala 92:32]
  wire  _T_642; // @[ROB.scala 68:36]
  wire  _T_643; // @[ROB.scala 68:20]
  wire  _T_644_valid; // @[ROB.scala 68:10]
  wire [3:0] _T_644_bits_addr; // @[ROB.scala 68:10]
  wire  _T_657; // @[ROB.scala 70:56]
  wire  _T_670; // @[ROB.scala 74:39]
  wire  _T_682; // @[ROB.scala 82:60]
  wire  _T_683; // @[ROB.scala 82:38]
  wire  _GEN_1262; // @[ROB.scala 98:31]
  wire  _GEN_1263; // @[ROB.scala 98:31]
  wire  _GEN_1264; // @[ROB.scala 94:29]
  wire  _GEN_1279; // @[ROB.scala 94:29]
  wire  _GEN_1280; // @[ROB.scala 92:32]
  wire  _T_686; // @[ROB.scala 106:15]
  wire [19:0] _GEN_1570; // @[ROB.scala 106:33]
  wire [4:0] _T_689; // @[ROB.scala 118:46]
  wire  _T_691; // @[ROB.scala 121:9]
  wire  _T_692; // @[ROB.scala 121:9]
  assign _T_3 = {{1'd0}, uncommited}; // @[ROB.scala 44:48]
  assign _T_4 = _T_3[3:0]; // @[ROB.scala 44:48]
  assign _GEN_16 = 4'h1 == _T_4 ? buf_1_data : buf_0_data; // @[ROB.scala 43:50]
  assign _GEN_20 = 4'h1 == _T_4 ? buf_1_inst_info_rd_addr : buf_0_inst_info_rd_addr; // @[ROB.scala 43:50]
  assign _GEN_25 = 4'h1 == _T_4 ? buf_1_inst_info_ctrl_rf_w : buf_0_inst_info_ctrl_rf_w; // @[ROB.scala 43:50]
  assign _GEN_31 = 4'h1 == _T_4 ? buf_1_committable : buf_0_committable; // @[ROB.scala 43:50]
  assign _GEN_32 = 4'h2 == _T_4 ? buf_2_data : _GEN_16; // @[ROB.scala 43:50]
  assign _GEN_36 = 4'h2 == _T_4 ? buf_2_inst_info_rd_addr : _GEN_20; // @[ROB.scala 43:50]
  assign _GEN_41 = 4'h2 == _T_4 ? buf_2_inst_info_ctrl_rf_w : _GEN_25; // @[ROB.scala 43:50]
  assign _GEN_47 = 4'h2 == _T_4 ? buf_2_committable : _GEN_31; // @[ROB.scala 43:50]
  assign _GEN_48 = 4'h3 == _T_4 ? buf_3_data : _GEN_32; // @[ROB.scala 43:50]
  assign _GEN_52 = 4'h3 == _T_4 ? buf_3_inst_info_rd_addr : _GEN_36; // @[ROB.scala 43:50]
  assign _GEN_57 = 4'h3 == _T_4 ? buf_3_inst_info_ctrl_rf_w : _GEN_41; // @[ROB.scala 43:50]
  assign _GEN_63 = 4'h3 == _T_4 ? buf_3_committable : _GEN_47; // @[ROB.scala 43:50]
  assign _GEN_64 = 4'h4 == _T_4 ? buf_4_data : _GEN_48; // @[ROB.scala 43:50]
  assign _GEN_68 = 4'h4 == _T_4 ? buf_4_inst_info_rd_addr : _GEN_52; // @[ROB.scala 43:50]
  assign _GEN_73 = 4'h4 == _T_4 ? buf_4_inst_info_ctrl_rf_w : _GEN_57; // @[ROB.scala 43:50]
  assign _GEN_79 = 4'h4 == _T_4 ? buf_4_committable : _GEN_63; // @[ROB.scala 43:50]
  assign _GEN_80 = 4'h5 == _T_4 ? buf_5_data : _GEN_64; // @[ROB.scala 43:50]
  assign _GEN_84 = 4'h5 == _T_4 ? buf_5_inst_info_rd_addr : _GEN_68; // @[ROB.scala 43:50]
  assign _GEN_89 = 4'h5 == _T_4 ? buf_5_inst_info_ctrl_rf_w : _GEN_73; // @[ROB.scala 43:50]
  assign _GEN_95 = 4'h5 == _T_4 ? buf_5_committable : _GEN_79; // @[ROB.scala 43:50]
  assign _GEN_96 = 4'h6 == _T_4 ? buf_6_data : _GEN_80; // @[ROB.scala 43:50]
  assign _GEN_100 = 4'h6 == _T_4 ? buf_6_inst_info_rd_addr : _GEN_84; // @[ROB.scala 43:50]
  assign _GEN_105 = 4'h6 == _T_4 ? buf_6_inst_info_ctrl_rf_w : _GEN_89; // @[ROB.scala 43:50]
  assign _GEN_111 = 4'h6 == _T_4 ? buf_6_committable : _GEN_95; // @[ROB.scala 43:50]
  assign _GEN_112 = 4'h7 == _T_4 ? buf_7_data : _GEN_96; // @[ROB.scala 43:50]
  assign _GEN_116 = 4'h7 == _T_4 ? buf_7_inst_info_rd_addr : _GEN_100; // @[ROB.scala 43:50]
  assign _GEN_121 = 4'h7 == _T_4 ? buf_7_inst_info_ctrl_rf_w : _GEN_105; // @[ROB.scala 43:50]
  assign _GEN_127 = 4'h7 == _T_4 ? buf_7_committable : _GEN_111; // @[ROB.scala 43:50]
  assign _GEN_128 = 4'h8 == _T_4 ? buf_8_data : _GEN_112; // @[ROB.scala 43:50]
  assign _GEN_132 = 4'h8 == _T_4 ? buf_8_inst_info_rd_addr : _GEN_116; // @[ROB.scala 43:50]
  assign _GEN_137 = 4'h8 == _T_4 ? buf_8_inst_info_ctrl_rf_w : _GEN_121; // @[ROB.scala 43:50]
  assign _GEN_143 = 4'h8 == _T_4 ? buf_8_committable : _GEN_127; // @[ROB.scala 43:50]
  assign _GEN_144 = 4'h9 == _T_4 ? buf_9_data : _GEN_128; // @[ROB.scala 43:50]
  assign _GEN_148 = 4'h9 == _T_4 ? buf_9_inst_info_rd_addr : _GEN_132; // @[ROB.scala 43:50]
  assign _GEN_153 = 4'h9 == _T_4 ? buf_9_inst_info_ctrl_rf_w : _GEN_137; // @[ROB.scala 43:50]
  assign _GEN_159 = 4'h9 == _T_4 ? buf_9_committable : _GEN_143; // @[ROB.scala 43:50]
  assign _GEN_160 = 4'ha == _T_4 ? buf_10_data : _GEN_144; // @[ROB.scala 43:50]
  assign _GEN_164 = 4'ha == _T_4 ? buf_10_inst_info_rd_addr : _GEN_148; // @[ROB.scala 43:50]
  assign _GEN_169 = 4'ha == _T_4 ? buf_10_inst_info_ctrl_rf_w : _GEN_153; // @[ROB.scala 43:50]
  assign _GEN_175 = 4'ha == _T_4 ? buf_10_committable : _GEN_159; // @[ROB.scala 43:50]
  assign _GEN_176 = 4'hb == _T_4 ? buf_11_data : _GEN_160; // @[ROB.scala 43:50]
  assign _GEN_180 = 4'hb == _T_4 ? buf_11_inst_info_rd_addr : _GEN_164; // @[ROB.scala 43:50]
  assign _GEN_185 = 4'hb == _T_4 ? buf_11_inst_info_ctrl_rf_w : _GEN_169; // @[ROB.scala 43:50]
  assign _GEN_191 = 4'hb == _T_4 ? buf_11_committable : _GEN_175; // @[ROB.scala 43:50]
  assign _GEN_192 = 4'hc == _T_4 ? buf_12_data : _GEN_176; // @[ROB.scala 43:50]
  assign _GEN_196 = 4'hc == _T_4 ? buf_12_inst_info_rd_addr : _GEN_180; // @[ROB.scala 43:50]
  assign _GEN_201 = 4'hc == _T_4 ? buf_12_inst_info_ctrl_rf_w : _GEN_185; // @[ROB.scala 43:50]
  assign _GEN_207 = 4'hc == _T_4 ? buf_12_committable : _GEN_191; // @[ROB.scala 43:50]
  assign _GEN_208 = 4'hd == _T_4 ? buf_13_data : _GEN_192; // @[ROB.scala 43:50]
  assign _GEN_212 = 4'hd == _T_4 ? buf_13_inst_info_rd_addr : _GEN_196; // @[ROB.scala 43:50]
  assign _GEN_217 = 4'hd == _T_4 ? buf_13_inst_info_ctrl_rf_w : _GEN_201; // @[ROB.scala 43:50]
  assign _GEN_223 = 4'hd == _T_4 ? buf_13_committable : _GEN_207; // @[ROB.scala 43:50]
  assign _GEN_224 = 4'he == _T_4 ? buf_14_data : _GEN_208; // @[ROB.scala 43:50]
  assign _GEN_228 = 4'he == _T_4 ? buf_14_inst_info_rd_addr : _GEN_212; // @[ROB.scala 43:50]
  assign _GEN_233 = 4'he == _T_4 ? buf_14_inst_info_ctrl_rf_w : _GEN_217; // @[ROB.scala 43:50]
  assign _GEN_239 = 4'he == _T_4 ? buf_14_committable : _GEN_223; // @[ROB.scala 43:50]
  assign _GEN_240 = 4'hf == _T_4 ? buf_15_data : _GEN_224; // @[ROB.scala 43:50]
  assign _GEN_244 = 4'hf == _T_4 ? buf_15_inst_info_rd_addr : _GEN_228; // @[ROB.scala 43:50]
  assign _GEN_249 = 4'hf == _T_4 ? buf_15_inst_info_ctrl_rf_w : _GEN_233; // @[ROB.scala 43:50]
  assign commitable_0 = 4'hf == _T_4 ? buf_15_committable : _GEN_239; // @[ROB.scala 43:50]
  assign _GEN_1571 = {{3'd0}, commitable_0}; // @[ROB.scala 50:41]
  assign next_uncommited = uncommited + _GEN_1571; // @[ROB.scala 50:41]
  assign _T_7 = io_graduate_0_valid & io_graduate_0_bits_mispredicted; // @[ROB.scala 53:136]
  assign _T_8_valid = _T_7 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 53:126]
  assign _T_8_bits_addr = _T_7 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 53:126]
  assign _T_8_bits_mispredicted = _T_7 & io_graduate_0_bits_mispredicted; // @[ROB.scala 53:126]
  assign mispredicted = _T_8_valid & _T_8_bits_mispredicted; // @[ROB.scala 54:53]
  assign _GEN_1572 = {{3'd0}, io_used_num}; // @[ROB.scala 58:46]
  assign unreserved_add_used = unreserved + _GEN_1572; // @[ROB.scala 58:46]
  assign _GEN_286 = 4'h1 == unreserved_add_used ? buf_1_reserved : buf_0_reserved; // @[ROB.scala 59:41]
  assign _GEN_302 = 4'h2 == unreserved_add_used ? buf_2_reserved : _GEN_286; // @[ROB.scala 59:41]
  assign _GEN_318 = 4'h3 == unreserved_add_used ? buf_3_reserved : _GEN_302; // @[ROB.scala 59:41]
  assign _GEN_334 = 4'h4 == unreserved_add_used ? buf_4_reserved : _GEN_318; // @[ROB.scala 59:41]
  assign _GEN_350 = 4'h5 == unreserved_add_used ? buf_5_reserved : _GEN_334; // @[ROB.scala 59:41]
  assign _GEN_366 = 4'h6 == unreserved_add_used ? buf_6_reserved : _GEN_350; // @[ROB.scala 59:41]
  assign _GEN_382 = 4'h7 == unreserved_add_used ? buf_7_reserved : _GEN_366; // @[ROB.scala 59:41]
  assign _GEN_398 = 4'h8 == unreserved_add_used ? buf_8_reserved : _GEN_382; // @[ROB.scala 59:41]
  assign _GEN_414 = 4'h9 == unreserved_add_used ? buf_9_reserved : _GEN_398; // @[ROB.scala 59:41]
  assign _GEN_430 = 4'ha == unreserved_add_used ? buf_10_reserved : _GEN_414; // @[ROB.scala 59:41]
  assign _GEN_446 = 4'hb == unreserved_add_used ? buf_11_reserved : _GEN_430; // @[ROB.scala 59:41]
  assign _GEN_462 = 4'hc == unreserved_add_used ? buf_12_reserved : _GEN_446; // @[ROB.scala 59:41]
  assign _GEN_478 = 4'hd == unreserved_add_used ? buf_13_reserved : _GEN_462; // @[ROB.scala 59:41]
  assign _GEN_494 = 4'he == unreserved_add_used ? buf_14_reserved : _GEN_478; // @[ROB.scala 59:41]
  assign _GEN_510 = 4'hf == unreserved_add_used ? buf_15_reserved : _GEN_494; // @[ROB.scala 59:41]
  assign unreserved_add_used_valid = _GEN_510 == 1'h0; // @[ROB.scala 59:41]
  assign _T_11 = unreserved_add_used_valid ? unreserved_add_used : unreserved; // @[Mux.scala 87:16]
  assign next_unreserved = mispredicted ? _T_8_bits_addr : _T_11; // @[Mux.scala 87:16]
  assign _T_12 = io_graduate_0_bits_addr == 4'h0; // @[ROB.scala 68:36]
  assign _T_13 = io_graduate_0_valid & _T_12; // @[ROB.scala 68:20]
  assign _T_14_valid = _T_13 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_14_bits_addr = _T_13 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_16 = _T_8_bits_addr <= unreserved; // @[ROB.scala 71:27]
  assign _T_17 = _T_8_bits_addr <= 4'h0; // @[ROB.scala 71:61]
  assign _T_18 = _T_16 & _T_17; // @[ROB.scala 71:41]
  assign _T_19 = 4'h0 < unreserved; // @[ROB.scala 71:75]
  assign _T_20 = _T_18 & _T_19; // @[ROB.scala 71:68]
  assign _T_21 = _T_8_bits_addr > unreserved; // @[ROB.scala 72:27]
  assign _T_24 = _T_19 | _T_17; // @[ROB.scala 72:61]
  assign _T_25 = _T_21 & _T_24; // @[ROB.scala 72:40]
  assign _T_26 = _T_20 | _T_25; // @[ROB.scala 71:89]
  assign _T_27 = mispredicted & _T_26; // @[ROB.scala 70:56]
  assign _T_28 = mispredicted == 1'h0; // @[ROB.scala 74:25]
  assign _T_29 = unreserved <= next_unreserved; // @[ROB.scala 75:20]
  assign _T_30 = unreserved <= 4'h0; // @[ROB.scala 75:55]
  assign _T_31 = 4'h0 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_32 = _T_30 & _T_31; // @[ROB.scala 75:62]
  assign _T_33 = _T_29 & _T_32; // @[ROB.scala 75:40]
  assign _T_34 = unreserved > next_unreserved; // @[ROB.scala 76:20]
  assign _T_37 = _T_31 | _T_30; // @[ROB.scala 76:65]
  assign _T_38 = _T_34 & _T_37; // @[ROB.scala 76:39]
  assign _T_39 = _T_33 | _T_38; // @[ROB.scala 75:89]
  assign _T_40 = _T_28 & _T_39; // @[ROB.scala 74:39]
  assign _T_41 = uncommited <= next_uncommited; // @[ROB.scala 79:20]
  assign _T_42 = uncommited <= 4'h0; // @[ROB.scala 79:55]
  assign _T_43 = 4'h0 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_44 = _T_42 & _T_43; // @[ROB.scala 79:62]
  assign _T_45 = _T_41 & _T_44; // @[ROB.scala 79:40]
  assign _T_46 = uncommited > next_uncommited; // @[ROB.scala 80:20]
  assign _T_49 = _T_43 | _T_42; // @[ROB.scala 80:66]
  assign _T_50 = _T_46 & _T_49; // @[ROB.scala 80:40]
  assign _T_51 = _T_45 | _T_50; // @[ROB.scala 79:89]
  assign _T_52 = _T_14_bits_addr == 4'h0; // @[ROB.scala 82:60]
  assign _T_53 = _T_14_valid & _T_52; // @[ROB.scala 82:38]
  assign _GEN_512 = _T_51 ? 1'h0 : buf_0_reserved; // @[ROB.scala 98:31]
  assign _GEN_513 = _T_51 ? 1'h0 : buf_0_committable; // @[ROB.scala 98:31]
  assign _GEN_514 = _T_53 | _GEN_513; // @[ROB.scala 94:29]
  assign _GEN_529 = _T_53 ? buf_0_reserved : _GEN_512; // @[ROB.scala 94:29]
  assign _GEN_530 = _T_40 | _GEN_529; // @[ROB.scala 92:32]
  assign _T_54 = io_graduate_0_bits_addr == 4'h1; // @[ROB.scala 68:36]
  assign _T_55 = io_graduate_0_valid & _T_54; // @[ROB.scala 68:20]
  assign _T_56_valid = _T_55 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_56_bits_addr = _T_55 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_59 = _T_8_bits_addr <= 4'h1; // @[ROB.scala 71:61]
  assign _T_60 = _T_16 & _T_59; // @[ROB.scala 71:41]
  assign _T_61 = 4'h1 < unreserved; // @[ROB.scala 71:75]
  assign _T_62 = _T_60 & _T_61; // @[ROB.scala 71:68]
  assign _T_66 = _T_61 | _T_59; // @[ROB.scala 72:61]
  assign _T_67 = _T_21 & _T_66; // @[ROB.scala 72:40]
  assign _T_68 = _T_62 | _T_67; // @[ROB.scala 71:89]
  assign _T_69 = mispredicted & _T_68; // @[ROB.scala 70:56]
  assign _T_72 = unreserved <= 4'h1; // @[ROB.scala 75:55]
  assign _T_73 = 4'h1 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_74 = _T_72 & _T_73; // @[ROB.scala 75:62]
  assign _T_75 = _T_29 & _T_74; // @[ROB.scala 75:40]
  assign _T_79 = _T_73 | _T_72; // @[ROB.scala 76:65]
  assign _T_80 = _T_34 & _T_79; // @[ROB.scala 76:39]
  assign _T_81 = _T_75 | _T_80; // @[ROB.scala 75:89]
  assign _T_82 = _T_28 & _T_81; // @[ROB.scala 74:39]
  assign _T_84 = uncommited <= 4'h1; // @[ROB.scala 79:55]
  assign _T_85 = 4'h1 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_86 = _T_84 & _T_85; // @[ROB.scala 79:62]
  assign _T_87 = _T_41 & _T_86; // @[ROB.scala 79:40]
  assign _T_91 = _T_85 | _T_84; // @[ROB.scala 80:66]
  assign _T_92 = _T_46 & _T_91; // @[ROB.scala 80:40]
  assign _T_93 = _T_87 | _T_92; // @[ROB.scala 79:89]
  assign _T_94 = _T_56_bits_addr == 4'h1; // @[ROB.scala 82:60]
  assign _T_95 = _T_56_valid & _T_94; // @[ROB.scala 82:38]
  assign _GEN_562 = _T_93 ? 1'h0 : buf_1_reserved; // @[ROB.scala 98:31]
  assign _GEN_563 = _T_93 ? 1'h0 : buf_1_committable; // @[ROB.scala 98:31]
  assign _GEN_564 = _T_95 | _GEN_563; // @[ROB.scala 94:29]
  assign _GEN_579 = _T_95 ? buf_1_reserved : _GEN_562; // @[ROB.scala 94:29]
  assign _GEN_580 = _T_82 | _GEN_579; // @[ROB.scala 92:32]
  assign _T_96 = io_graduate_0_bits_addr == 4'h2; // @[ROB.scala 68:36]
  assign _T_97 = io_graduate_0_valid & _T_96; // @[ROB.scala 68:20]
  assign _T_98_valid = _T_97 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_98_bits_addr = _T_97 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_101 = _T_8_bits_addr <= 4'h2; // @[ROB.scala 71:61]
  assign _T_102 = _T_16 & _T_101; // @[ROB.scala 71:41]
  assign _T_103 = 4'h2 < unreserved; // @[ROB.scala 71:75]
  assign _T_104 = _T_102 & _T_103; // @[ROB.scala 71:68]
  assign _T_108 = _T_103 | _T_101; // @[ROB.scala 72:61]
  assign _T_109 = _T_21 & _T_108; // @[ROB.scala 72:40]
  assign _T_110 = _T_104 | _T_109; // @[ROB.scala 71:89]
  assign _T_111 = mispredicted & _T_110; // @[ROB.scala 70:56]
  assign _T_114 = unreserved <= 4'h2; // @[ROB.scala 75:55]
  assign _T_115 = 4'h2 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_116 = _T_114 & _T_115; // @[ROB.scala 75:62]
  assign _T_117 = _T_29 & _T_116; // @[ROB.scala 75:40]
  assign _T_121 = _T_115 | _T_114; // @[ROB.scala 76:65]
  assign _T_122 = _T_34 & _T_121; // @[ROB.scala 76:39]
  assign _T_123 = _T_117 | _T_122; // @[ROB.scala 75:89]
  assign _T_124 = _T_28 & _T_123; // @[ROB.scala 74:39]
  assign _T_126 = uncommited <= 4'h2; // @[ROB.scala 79:55]
  assign _T_127 = 4'h2 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_128 = _T_126 & _T_127; // @[ROB.scala 79:62]
  assign _T_129 = _T_41 & _T_128; // @[ROB.scala 79:40]
  assign _T_133 = _T_127 | _T_126; // @[ROB.scala 80:66]
  assign _T_134 = _T_46 & _T_133; // @[ROB.scala 80:40]
  assign _T_135 = _T_129 | _T_134; // @[ROB.scala 79:89]
  assign _T_136 = _T_98_bits_addr == 4'h2; // @[ROB.scala 82:60]
  assign _T_137 = _T_98_valid & _T_136; // @[ROB.scala 82:38]
  assign _GEN_612 = _T_135 ? 1'h0 : buf_2_reserved; // @[ROB.scala 98:31]
  assign _GEN_613 = _T_135 ? 1'h0 : buf_2_committable; // @[ROB.scala 98:31]
  assign _GEN_614 = _T_137 | _GEN_613; // @[ROB.scala 94:29]
  assign _GEN_629 = _T_137 ? buf_2_reserved : _GEN_612; // @[ROB.scala 94:29]
  assign _GEN_630 = _T_124 | _GEN_629; // @[ROB.scala 92:32]
  assign _T_138 = io_graduate_0_bits_addr == 4'h3; // @[ROB.scala 68:36]
  assign _T_139 = io_graduate_0_valid & _T_138; // @[ROB.scala 68:20]
  assign _T_140_valid = _T_139 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_140_bits_addr = _T_139 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_143 = _T_8_bits_addr <= 4'h3; // @[ROB.scala 71:61]
  assign _T_144 = _T_16 & _T_143; // @[ROB.scala 71:41]
  assign _T_145 = 4'h3 < unreserved; // @[ROB.scala 71:75]
  assign _T_146 = _T_144 & _T_145; // @[ROB.scala 71:68]
  assign _T_150 = _T_145 | _T_143; // @[ROB.scala 72:61]
  assign _T_151 = _T_21 & _T_150; // @[ROB.scala 72:40]
  assign _T_152 = _T_146 | _T_151; // @[ROB.scala 71:89]
  assign _T_153 = mispredicted & _T_152; // @[ROB.scala 70:56]
  assign _T_156 = unreserved <= 4'h3; // @[ROB.scala 75:55]
  assign _T_157 = 4'h3 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_158 = _T_156 & _T_157; // @[ROB.scala 75:62]
  assign _T_159 = _T_29 & _T_158; // @[ROB.scala 75:40]
  assign _T_163 = _T_157 | _T_156; // @[ROB.scala 76:65]
  assign _T_164 = _T_34 & _T_163; // @[ROB.scala 76:39]
  assign _T_165 = _T_159 | _T_164; // @[ROB.scala 75:89]
  assign _T_166 = _T_28 & _T_165; // @[ROB.scala 74:39]
  assign _T_168 = uncommited <= 4'h3; // @[ROB.scala 79:55]
  assign _T_169 = 4'h3 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_170 = _T_168 & _T_169; // @[ROB.scala 79:62]
  assign _T_171 = _T_41 & _T_170; // @[ROB.scala 79:40]
  assign _T_175 = _T_169 | _T_168; // @[ROB.scala 80:66]
  assign _T_176 = _T_46 & _T_175; // @[ROB.scala 80:40]
  assign _T_177 = _T_171 | _T_176; // @[ROB.scala 79:89]
  assign _T_178 = _T_140_bits_addr == 4'h3; // @[ROB.scala 82:60]
  assign _T_179 = _T_140_valid & _T_178; // @[ROB.scala 82:38]
  assign _GEN_662 = _T_177 ? 1'h0 : buf_3_reserved; // @[ROB.scala 98:31]
  assign _GEN_663 = _T_177 ? 1'h0 : buf_3_committable; // @[ROB.scala 98:31]
  assign _GEN_664 = _T_179 | _GEN_663; // @[ROB.scala 94:29]
  assign _GEN_679 = _T_179 ? buf_3_reserved : _GEN_662; // @[ROB.scala 94:29]
  assign _GEN_680 = _T_166 | _GEN_679; // @[ROB.scala 92:32]
  assign _T_180 = io_graduate_0_bits_addr == 4'h4; // @[ROB.scala 68:36]
  assign _T_181 = io_graduate_0_valid & _T_180; // @[ROB.scala 68:20]
  assign _T_182_valid = _T_181 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_182_bits_addr = _T_181 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_185 = _T_8_bits_addr <= 4'h4; // @[ROB.scala 71:61]
  assign _T_186 = _T_16 & _T_185; // @[ROB.scala 71:41]
  assign _T_187 = 4'h4 < unreserved; // @[ROB.scala 71:75]
  assign _T_188 = _T_186 & _T_187; // @[ROB.scala 71:68]
  assign _T_192 = _T_187 | _T_185; // @[ROB.scala 72:61]
  assign _T_193 = _T_21 & _T_192; // @[ROB.scala 72:40]
  assign _T_194 = _T_188 | _T_193; // @[ROB.scala 71:89]
  assign _T_195 = mispredicted & _T_194; // @[ROB.scala 70:56]
  assign _T_198 = unreserved <= 4'h4; // @[ROB.scala 75:55]
  assign _T_199 = 4'h4 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_200 = _T_198 & _T_199; // @[ROB.scala 75:62]
  assign _T_201 = _T_29 & _T_200; // @[ROB.scala 75:40]
  assign _T_205 = _T_199 | _T_198; // @[ROB.scala 76:65]
  assign _T_206 = _T_34 & _T_205; // @[ROB.scala 76:39]
  assign _T_207 = _T_201 | _T_206; // @[ROB.scala 75:89]
  assign _T_208 = _T_28 & _T_207; // @[ROB.scala 74:39]
  assign _T_210 = uncommited <= 4'h4; // @[ROB.scala 79:55]
  assign _T_211 = 4'h4 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_212 = _T_210 & _T_211; // @[ROB.scala 79:62]
  assign _T_213 = _T_41 & _T_212; // @[ROB.scala 79:40]
  assign _T_217 = _T_211 | _T_210; // @[ROB.scala 80:66]
  assign _T_218 = _T_46 & _T_217; // @[ROB.scala 80:40]
  assign _T_219 = _T_213 | _T_218; // @[ROB.scala 79:89]
  assign _T_220 = _T_182_bits_addr == 4'h4; // @[ROB.scala 82:60]
  assign _T_221 = _T_182_valid & _T_220; // @[ROB.scala 82:38]
  assign _GEN_712 = _T_219 ? 1'h0 : buf_4_reserved; // @[ROB.scala 98:31]
  assign _GEN_713 = _T_219 ? 1'h0 : buf_4_committable; // @[ROB.scala 98:31]
  assign _GEN_714 = _T_221 | _GEN_713; // @[ROB.scala 94:29]
  assign _GEN_729 = _T_221 ? buf_4_reserved : _GEN_712; // @[ROB.scala 94:29]
  assign _GEN_730 = _T_208 | _GEN_729; // @[ROB.scala 92:32]
  assign _T_222 = io_graduate_0_bits_addr == 4'h5; // @[ROB.scala 68:36]
  assign _T_223 = io_graduate_0_valid & _T_222; // @[ROB.scala 68:20]
  assign _T_224_valid = _T_223 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_224_bits_addr = _T_223 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_227 = _T_8_bits_addr <= 4'h5; // @[ROB.scala 71:61]
  assign _T_228 = _T_16 & _T_227; // @[ROB.scala 71:41]
  assign _T_229 = 4'h5 < unreserved; // @[ROB.scala 71:75]
  assign _T_230 = _T_228 & _T_229; // @[ROB.scala 71:68]
  assign _T_234 = _T_229 | _T_227; // @[ROB.scala 72:61]
  assign _T_235 = _T_21 & _T_234; // @[ROB.scala 72:40]
  assign _T_236 = _T_230 | _T_235; // @[ROB.scala 71:89]
  assign _T_237 = mispredicted & _T_236; // @[ROB.scala 70:56]
  assign _T_240 = unreserved <= 4'h5; // @[ROB.scala 75:55]
  assign _T_241 = 4'h5 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_242 = _T_240 & _T_241; // @[ROB.scala 75:62]
  assign _T_243 = _T_29 & _T_242; // @[ROB.scala 75:40]
  assign _T_247 = _T_241 | _T_240; // @[ROB.scala 76:65]
  assign _T_248 = _T_34 & _T_247; // @[ROB.scala 76:39]
  assign _T_249 = _T_243 | _T_248; // @[ROB.scala 75:89]
  assign _T_250 = _T_28 & _T_249; // @[ROB.scala 74:39]
  assign _T_252 = uncommited <= 4'h5; // @[ROB.scala 79:55]
  assign _T_253 = 4'h5 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_254 = _T_252 & _T_253; // @[ROB.scala 79:62]
  assign _T_255 = _T_41 & _T_254; // @[ROB.scala 79:40]
  assign _T_259 = _T_253 | _T_252; // @[ROB.scala 80:66]
  assign _T_260 = _T_46 & _T_259; // @[ROB.scala 80:40]
  assign _T_261 = _T_255 | _T_260; // @[ROB.scala 79:89]
  assign _T_262 = _T_224_bits_addr == 4'h5; // @[ROB.scala 82:60]
  assign _T_263 = _T_224_valid & _T_262; // @[ROB.scala 82:38]
  assign _GEN_762 = _T_261 ? 1'h0 : buf_5_reserved; // @[ROB.scala 98:31]
  assign _GEN_763 = _T_261 ? 1'h0 : buf_5_committable; // @[ROB.scala 98:31]
  assign _GEN_764 = _T_263 | _GEN_763; // @[ROB.scala 94:29]
  assign _GEN_779 = _T_263 ? buf_5_reserved : _GEN_762; // @[ROB.scala 94:29]
  assign _GEN_780 = _T_250 | _GEN_779; // @[ROB.scala 92:32]
  assign _T_264 = io_graduate_0_bits_addr == 4'h6; // @[ROB.scala 68:36]
  assign _T_265 = io_graduate_0_valid & _T_264; // @[ROB.scala 68:20]
  assign _T_266_valid = _T_265 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_266_bits_addr = _T_265 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_269 = _T_8_bits_addr <= 4'h6; // @[ROB.scala 71:61]
  assign _T_270 = _T_16 & _T_269; // @[ROB.scala 71:41]
  assign _T_271 = 4'h6 < unreserved; // @[ROB.scala 71:75]
  assign _T_272 = _T_270 & _T_271; // @[ROB.scala 71:68]
  assign _T_276 = _T_271 | _T_269; // @[ROB.scala 72:61]
  assign _T_277 = _T_21 & _T_276; // @[ROB.scala 72:40]
  assign _T_278 = _T_272 | _T_277; // @[ROB.scala 71:89]
  assign _T_279 = mispredicted & _T_278; // @[ROB.scala 70:56]
  assign _T_282 = unreserved <= 4'h6; // @[ROB.scala 75:55]
  assign _T_283 = 4'h6 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_284 = _T_282 & _T_283; // @[ROB.scala 75:62]
  assign _T_285 = _T_29 & _T_284; // @[ROB.scala 75:40]
  assign _T_289 = _T_283 | _T_282; // @[ROB.scala 76:65]
  assign _T_290 = _T_34 & _T_289; // @[ROB.scala 76:39]
  assign _T_291 = _T_285 | _T_290; // @[ROB.scala 75:89]
  assign _T_292 = _T_28 & _T_291; // @[ROB.scala 74:39]
  assign _T_294 = uncommited <= 4'h6; // @[ROB.scala 79:55]
  assign _T_295 = 4'h6 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_296 = _T_294 & _T_295; // @[ROB.scala 79:62]
  assign _T_297 = _T_41 & _T_296; // @[ROB.scala 79:40]
  assign _T_301 = _T_295 | _T_294; // @[ROB.scala 80:66]
  assign _T_302 = _T_46 & _T_301; // @[ROB.scala 80:40]
  assign _T_303 = _T_297 | _T_302; // @[ROB.scala 79:89]
  assign _T_304 = _T_266_bits_addr == 4'h6; // @[ROB.scala 82:60]
  assign _T_305 = _T_266_valid & _T_304; // @[ROB.scala 82:38]
  assign _GEN_812 = _T_303 ? 1'h0 : buf_6_reserved; // @[ROB.scala 98:31]
  assign _GEN_813 = _T_303 ? 1'h0 : buf_6_committable; // @[ROB.scala 98:31]
  assign _GEN_814 = _T_305 | _GEN_813; // @[ROB.scala 94:29]
  assign _GEN_829 = _T_305 ? buf_6_reserved : _GEN_812; // @[ROB.scala 94:29]
  assign _GEN_830 = _T_292 | _GEN_829; // @[ROB.scala 92:32]
  assign _T_306 = io_graduate_0_bits_addr == 4'h7; // @[ROB.scala 68:36]
  assign _T_307 = io_graduate_0_valid & _T_306; // @[ROB.scala 68:20]
  assign _T_308_valid = _T_307 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_308_bits_addr = _T_307 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_311 = _T_8_bits_addr <= 4'h7; // @[ROB.scala 71:61]
  assign _T_312 = _T_16 & _T_311; // @[ROB.scala 71:41]
  assign _T_313 = 4'h7 < unreserved; // @[ROB.scala 71:75]
  assign _T_314 = _T_312 & _T_313; // @[ROB.scala 71:68]
  assign _T_318 = _T_313 | _T_311; // @[ROB.scala 72:61]
  assign _T_319 = _T_21 & _T_318; // @[ROB.scala 72:40]
  assign _T_320 = _T_314 | _T_319; // @[ROB.scala 71:89]
  assign _T_321 = mispredicted & _T_320; // @[ROB.scala 70:56]
  assign _T_324 = unreserved <= 4'h7; // @[ROB.scala 75:55]
  assign _T_325 = 4'h7 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_326 = _T_324 & _T_325; // @[ROB.scala 75:62]
  assign _T_327 = _T_29 & _T_326; // @[ROB.scala 75:40]
  assign _T_331 = _T_325 | _T_324; // @[ROB.scala 76:65]
  assign _T_332 = _T_34 & _T_331; // @[ROB.scala 76:39]
  assign _T_333 = _T_327 | _T_332; // @[ROB.scala 75:89]
  assign _T_334 = _T_28 & _T_333; // @[ROB.scala 74:39]
  assign _T_336 = uncommited <= 4'h7; // @[ROB.scala 79:55]
  assign _T_337 = 4'h7 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_338 = _T_336 & _T_337; // @[ROB.scala 79:62]
  assign _T_339 = _T_41 & _T_338; // @[ROB.scala 79:40]
  assign _T_343 = _T_337 | _T_336; // @[ROB.scala 80:66]
  assign _T_344 = _T_46 & _T_343; // @[ROB.scala 80:40]
  assign _T_345 = _T_339 | _T_344; // @[ROB.scala 79:89]
  assign _T_346 = _T_308_bits_addr == 4'h7; // @[ROB.scala 82:60]
  assign _T_347 = _T_308_valid & _T_346; // @[ROB.scala 82:38]
  assign _GEN_862 = _T_345 ? 1'h0 : buf_7_reserved; // @[ROB.scala 98:31]
  assign _GEN_863 = _T_345 ? 1'h0 : buf_7_committable; // @[ROB.scala 98:31]
  assign _GEN_864 = _T_347 | _GEN_863; // @[ROB.scala 94:29]
  assign _GEN_879 = _T_347 ? buf_7_reserved : _GEN_862; // @[ROB.scala 94:29]
  assign _GEN_880 = _T_334 | _GEN_879; // @[ROB.scala 92:32]
  assign _T_348 = io_graduate_0_bits_addr == 4'h8; // @[ROB.scala 68:36]
  assign _T_349 = io_graduate_0_valid & _T_348; // @[ROB.scala 68:20]
  assign _T_350_valid = _T_349 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_350_bits_addr = _T_349 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_353 = _T_8_bits_addr <= 4'h8; // @[ROB.scala 71:61]
  assign _T_354 = _T_16 & _T_353; // @[ROB.scala 71:41]
  assign _T_355 = 4'h8 < unreserved; // @[ROB.scala 71:75]
  assign _T_356 = _T_354 & _T_355; // @[ROB.scala 71:68]
  assign _T_360 = _T_355 | _T_353; // @[ROB.scala 72:61]
  assign _T_361 = _T_21 & _T_360; // @[ROB.scala 72:40]
  assign _T_362 = _T_356 | _T_361; // @[ROB.scala 71:89]
  assign _T_363 = mispredicted & _T_362; // @[ROB.scala 70:56]
  assign _T_366 = unreserved <= 4'h8; // @[ROB.scala 75:55]
  assign _T_367 = 4'h8 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_368 = _T_366 & _T_367; // @[ROB.scala 75:62]
  assign _T_369 = _T_29 & _T_368; // @[ROB.scala 75:40]
  assign _T_373 = _T_367 | _T_366; // @[ROB.scala 76:65]
  assign _T_374 = _T_34 & _T_373; // @[ROB.scala 76:39]
  assign _T_375 = _T_369 | _T_374; // @[ROB.scala 75:89]
  assign _T_376 = _T_28 & _T_375; // @[ROB.scala 74:39]
  assign _T_378 = uncommited <= 4'h8; // @[ROB.scala 79:55]
  assign _T_379 = 4'h8 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_380 = _T_378 & _T_379; // @[ROB.scala 79:62]
  assign _T_381 = _T_41 & _T_380; // @[ROB.scala 79:40]
  assign _T_385 = _T_379 | _T_378; // @[ROB.scala 80:66]
  assign _T_386 = _T_46 & _T_385; // @[ROB.scala 80:40]
  assign _T_387 = _T_381 | _T_386; // @[ROB.scala 79:89]
  assign _T_388 = _T_350_bits_addr == 4'h8; // @[ROB.scala 82:60]
  assign _T_389 = _T_350_valid & _T_388; // @[ROB.scala 82:38]
  assign _GEN_912 = _T_387 ? 1'h0 : buf_8_reserved; // @[ROB.scala 98:31]
  assign _GEN_913 = _T_387 ? 1'h0 : buf_8_committable; // @[ROB.scala 98:31]
  assign _GEN_914 = _T_389 | _GEN_913; // @[ROB.scala 94:29]
  assign _GEN_929 = _T_389 ? buf_8_reserved : _GEN_912; // @[ROB.scala 94:29]
  assign _GEN_930 = _T_376 | _GEN_929; // @[ROB.scala 92:32]
  assign _T_390 = io_graduate_0_bits_addr == 4'h9; // @[ROB.scala 68:36]
  assign _T_391 = io_graduate_0_valid & _T_390; // @[ROB.scala 68:20]
  assign _T_392_valid = _T_391 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_392_bits_addr = _T_391 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_395 = _T_8_bits_addr <= 4'h9; // @[ROB.scala 71:61]
  assign _T_396 = _T_16 & _T_395; // @[ROB.scala 71:41]
  assign _T_397 = 4'h9 < unreserved; // @[ROB.scala 71:75]
  assign _T_398 = _T_396 & _T_397; // @[ROB.scala 71:68]
  assign _T_402 = _T_397 | _T_395; // @[ROB.scala 72:61]
  assign _T_403 = _T_21 & _T_402; // @[ROB.scala 72:40]
  assign _T_404 = _T_398 | _T_403; // @[ROB.scala 71:89]
  assign _T_405 = mispredicted & _T_404; // @[ROB.scala 70:56]
  assign _T_408 = unreserved <= 4'h9; // @[ROB.scala 75:55]
  assign _T_409 = 4'h9 < next_unreserved; // @[ROB.scala 75:69]
  assign _T_410 = _T_408 & _T_409; // @[ROB.scala 75:62]
  assign _T_411 = _T_29 & _T_410; // @[ROB.scala 75:40]
  assign _T_415 = _T_409 | _T_408; // @[ROB.scala 76:65]
  assign _T_416 = _T_34 & _T_415; // @[ROB.scala 76:39]
  assign _T_417 = _T_411 | _T_416; // @[ROB.scala 75:89]
  assign _T_418 = _T_28 & _T_417; // @[ROB.scala 74:39]
  assign _T_420 = uncommited <= 4'h9; // @[ROB.scala 79:55]
  assign _T_421 = 4'h9 < next_uncommited; // @[ROB.scala 79:69]
  assign _T_422 = _T_420 & _T_421; // @[ROB.scala 79:62]
  assign _T_423 = _T_41 & _T_422; // @[ROB.scala 79:40]
  assign _T_427 = _T_421 | _T_420; // @[ROB.scala 80:66]
  assign _T_428 = _T_46 & _T_427; // @[ROB.scala 80:40]
  assign _T_429 = _T_423 | _T_428; // @[ROB.scala 79:89]
  assign _T_430 = _T_392_bits_addr == 4'h9; // @[ROB.scala 82:60]
  assign _T_431 = _T_392_valid & _T_430; // @[ROB.scala 82:38]
  assign _GEN_962 = _T_429 ? 1'h0 : buf_9_reserved; // @[ROB.scala 98:31]
  assign _GEN_963 = _T_429 ? 1'h0 : buf_9_committable; // @[ROB.scala 98:31]
  assign _GEN_964 = _T_431 | _GEN_963; // @[ROB.scala 94:29]
  assign _GEN_979 = _T_431 ? buf_9_reserved : _GEN_962; // @[ROB.scala 94:29]
  assign _GEN_980 = _T_418 | _GEN_979; // @[ROB.scala 92:32]
  assign _T_432 = io_graduate_0_bits_addr == 4'ha; // @[ROB.scala 68:36]
  assign _T_433 = io_graduate_0_valid & _T_432; // @[ROB.scala 68:20]
  assign _T_434_valid = _T_433 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_434_bits_addr = _T_433 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_437 = _T_8_bits_addr <= 4'ha; // @[ROB.scala 71:61]
  assign _T_438 = _T_16 & _T_437; // @[ROB.scala 71:41]
  assign _T_439 = 4'ha < unreserved; // @[ROB.scala 71:75]
  assign _T_440 = _T_438 & _T_439; // @[ROB.scala 71:68]
  assign _T_444 = _T_439 | _T_437; // @[ROB.scala 72:61]
  assign _T_445 = _T_21 & _T_444; // @[ROB.scala 72:40]
  assign _T_446 = _T_440 | _T_445; // @[ROB.scala 71:89]
  assign _T_447 = mispredicted & _T_446; // @[ROB.scala 70:56]
  assign _T_450 = unreserved <= 4'ha; // @[ROB.scala 75:55]
  assign _T_451 = 4'ha < next_unreserved; // @[ROB.scala 75:69]
  assign _T_452 = _T_450 & _T_451; // @[ROB.scala 75:62]
  assign _T_453 = _T_29 & _T_452; // @[ROB.scala 75:40]
  assign _T_457 = _T_451 | _T_450; // @[ROB.scala 76:65]
  assign _T_458 = _T_34 & _T_457; // @[ROB.scala 76:39]
  assign _T_459 = _T_453 | _T_458; // @[ROB.scala 75:89]
  assign _T_460 = _T_28 & _T_459; // @[ROB.scala 74:39]
  assign _T_462 = uncommited <= 4'ha; // @[ROB.scala 79:55]
  assign _T_463 = 4'ha < next_uncommited; // @[ROB.scala 79:69]
  assign _T_464 = _T_462 & _T_463; // @[ROB.scala 79:62]
  assign _T_465 = _T_41 & _T_464; // @[ROB.scala 79:40]
  assign _T_469 = _T_463 | _T_462; // @[ROB.scala 80:66]
  assign _T_470 = _T_46 & _T_469; // @[ROB.scala 80:40]
  assign _T_471 = _T_465 | _T_470; // @[ROB.scala 79:89]
  assign _T_472 = _T_434_bits_addr == 4'ha; // @[ROB.scala 82:60]
  assign _T_473 = _T_434_valid & _T_472; // @[ROB.scala 82:38]
  assign _GEN_1012 = _T_471 ? 1'h0 : buf_10_reserved; // @[ROB.scala 98:31]
  assign _GEN_1013 = _T_471 ? 1'h0 : buf_10_committable; // @[ROB.scala 98:31]
  assign _GEN_1014 = _T_473 | _GEN_1013; // @[ROB.scala 94:29]
  assign _GEN_1029 = _T_473 ? buf_10_reserved : _GEN_1012; // @[ROB.scala 94:29]
  assign _GEN_1030 = _T_460 | _GEN_1029; // @[ROB.scala 92:32]
  assign _T_474 = io_graduate_0_bits_addr == 4'hb; // @[ROB.scala 68:36]
  assign _T_475 = io_graduate_0_valid & _T_474; // @[ROB.scala 68:20]
  assign _T_476_valid = _T_475 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_476_bits_addr = _T_475 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_479 = _T_8_bits_addr <= 4'hb; // @[ROB.scala 71:61]
  assign _T_480 = _T_16 & _T_479; // @[ROB.scala 71:41]
  assign _T_481 = 4'hb < unreserved; // @[ROB.scala 71:75]
  assign _T_482 = _T_480 & _T_481; // @[ROB.scala 71:68]
  assign _T_486 = _T_481 | _T_479; // @[ROB.scala 72:61]
  assign _T_487 = _T_21 & _T_486; // @[ROB.scala 72:40]
  assign _T_488 = _T_482 | _T_487; // @[ROB.scala 71:89]
  assign _T_489 = mispredicted & _T_488; // @[ROB.scala 70:56]
  assign _T_492 = unreserved <= 4'hb; // @[ROB.scala 75:55]
  assign _T_493 = 4'hb < next_unreserved; // @[ROB.scala 75:69]
  assign _T_494 = _T_492 & _T_493; // @[ROB.scala 75:62]
  assign _T_495 = _T_29 & _T_494; // @[ROB.scala 75:40]
  assign _T_499 = _T_493 | _T_492; // @[ROB.scala 76:65]
  assign _T_500 = _T_34 & _T_499; // @[ROB.scala 76:39]
  assign _T_501 = _T_495 | _T_500; // @[ROB.scala 75:89]
  assign _T_502 = _T_28 & _T_501; // @[ROB.scala 74:39]
  assign _T_504 = uncommited <= 4'hb; // @[ROB.scala 79:55]
  assign _T_505 = 4'hb < next_uncommited; // @[ROB.scala 79:69]
  assign _T_506 = _T_504 & _T_505; // @[ROB.scala 79:62]
  assign _T_507 = _T_41 & _T_506; // @[ROB.scala 79:40]
  assign _T_511 = _T_505 | _T_504; // @[ROB.scala 80:66]
  assign _T_512 = _T_46 & _T_511; // @[ROB.scala 80:40]
  assign _T_513 = _T_507 | _T_512; // @[ROB.scala 79:89]
  assign _T_514 = _T_476_bits_addr == 4'hb; // @[ROB.scala 82:60]
  assign _T_515 = _T_476_valid & _T_514; // @[ROB.scala 82:38]
  assign _GEN_1062 = _T_513 ? 1'h0 : buf_11_reserved; // @[ROB.scala 98:31]
  assign _GEN_1063 = _T_513 ? 1'h0 : buf_11_committable; // @[ROB.scala 98:31]
  assign _GEN_1064 = _T_515 | _GEN_1063; // @[ROB.scala 94:29]
  assign _GEN_1079 = _T_515 ? buf_11_reserved : _GEN_1062; // @[ROB.scala 94:29]
  assign _GEN_1080 = _T_502 | _GEN_1079; // @[ROB.scala 92:32]
  assign _T_516 = io_graduate_0_bits_addr == 4'hc; // @[ROB.scala 68:36]
  assign _T_517 = io_graduate_0_valid & _T_516; // @[ROB.scala 68:20]
  assign _T_518_valid = _T_517 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_518_bits_addr = _T_517 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_521 = _T_8_bits_addr <= 4'hc; // @[ROB.scala 71:61]
  assign _T_522 = _T_16 & _T_521; // @[ROB.scala 71:41]
  assign _T_523 = 4'hc < unreserved; // @[ROB.scala 71:75]
  assign _T_524 = _T_522 & _T_523; // @[ROB.scala 71:68]
  assign _T_528 = _T_523 | _T_521; // @[ROB.scala 72:61]
  assign _T_529 = _T_21 & _T_528; // @[ROB.scala 72:40]
  assign _T_530 = _T_524 | _T_529; // @[ROB.scala 71:89]
  assign _T_531 = mispredicted & _T_530; // @[ROB.scala 70:56]
  assign _T_534 = unreserved <= 4'hc; // @[ROB.scala 75:55]
  assign _T_535 = 4'hc < next_unreserved; // @[ROB.scala 75:69]
  assign _T_536 = _T_534 & _T_535; // @[ROB.scala 75:62]
  assign _T_537 = _T_29 & _T_536; // @[ROB.scala 75:40]
  assign _T_541 = _T_535 | _T_534; // @[ROB.scala 76:65]
  assign _T_542 = _T_34 & _T_541; // @[ROB.scala 76:39]
  assign _T_543 = _T_537 | _T_542; // @[ROB.scala 75:89]
  assign _T_544 = _T_28 & _T_543; // @[ROB.scala 74:39]
  assign _T_546 = uncommited <= 4'hc; // @[ROB.scala 79:55]
  assign _T_547 = 4'hc < next_uncommited; // @[ROB.scala 79:69]
  assign _T_548 = _T_546 & _T_547; // @[ROB.scala 79:62]
  assign _T_549 = _T_41 & _T_548; // @[ROB.scala 79:40]
  assign _T_553 = _T_547 | _T_546; // @[ROB.scala 80:66]
  assign _T_554 = _T_46 & _T_553; // @[ROB.scala 80:40]
  assign _T_555 = _T_549 | _T_554; // @[ROB.scala 79:89]
  assign _T_556 = _T_518_bits_addr == 4'hc; // @[ROB.scala 82:60]
  assign _T_557 = _T_518_valid & _T_556; // @[ROB.scala 82:38]
  assign _GEN_1112 = _T_555 ? 1'h0 : buf_12_reserved; // @[ROB.scala 98:31]
  assign _GEN_1113 = _T_555 ? 1'h0 : buf_12_committable; // @[ROB.scala 98:31]
  assign _GEN_1114 = _T_557 | _GEN_1113; // @[ROB.scala 94:29]
  assign _GEN_1129 = _T_557 ? buf_12_reserved : _GEN_1112; // @[ROB.scala 94:29]
  assign _GEN_1130 = _T_544 | _GEN_1129; // @[ROB.scala 92:32]
  assign _T_558 = io_graduate_0_bits_addr == 4'hd; // @[ROB.scala 68:36]
  assign _T_559 = io_graduate_0_valid & _T_558; // @[ROB.scala 68:20]
  assign _T_560_valid = _T_559 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_560_bits_addr = _T_559 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_563 = _T_8_bits_addr <= 4'hd; // @[ROB.scala 71:61]
  assign _T_564 = _T_16 & _T_563; // @[ROB.scala 71:41]
  assign _T_565 = 4'hd < unreserved; // @[ROB.scala 71:75]
  assign _T_566 = _T_564 & _T_565; // @[ROB.scala 71:68]
  assign _T_570 = _T_565 | _T_563; // @[ROB.scala 72:61]
  assign _T_571 = _T_21 & _T_570; // @[ROB.scala 72:40]
  assign _T_572 = _T_566 | _T_571; // @[ROB.scala 71:89]
  assign _T_573 = mispredicted & _T_572; // @[ROB.scala 70:56]
  assign _T_576 = unreserved <= 4'hd; // @[ROB.scala 75:55]
  assign _T_577 = 4'hd < next_unreserved; // @[ROB.scala 75:69]
  assign _T_578 = _T_576 & _T_577; // @[ROB.scala 75:62]
  assign _T_579 = _T_29 & _T_578; // @[ROB.scala 75:40]
  assign _T_583 = _T_577 | _T_576; // @[ROB.scala 76:65]
  assign _T_584 = _T_34 & _T_583; // @[ROB.scala 76:39]
  assign _T_585 = _T_579 | _T_584; // @[ROB.scala 75:89]
  assign _T_586 = _T_28 & _T_585; // @[ROB.scala 74:39]
  assign _T_588 = uncommited <= 4'hd; // @[ROB.scala 79:55]
  assign _T_589 = 4'hd < next_uncommited; // @[ROB.scala 79:69]
  assign _T_590 = _T_588 & _T_589; // @[ROB.scala 79:62]
  assign _T_591 = _T_41 & _T_590; // @[ROB.scala 79:40]
  assign _T_595 = _T_589 | _T_588; // @[ROB.scala 80:66]
  assign _T_596 = _T_46 & _T_595; // @[ROB.scala 80:40]
  assign _T_597 = _T_591 | _T_596; // @[ROB.scala 79:89]
  assign _T_598 = _T_560_bits_addr == 4'hd; // @[ROB.scala 82:60]
  assign _T_599 = _T_560_valid & _T_598; // @[ROB.scala 82:38]
  assign _GEN_1162 = _T_597 ? 1'h0 : buf_13_reserved; // @[ROB.scala 98:31]
  assign _GEN_1163 = _T_597 ? 1'h0 : buf_13_committable; // @[ROB.scala 98:31]
  assign _GEN_1164 = _T_599 | _GEN_1163; // @[ROB.scala 94:29]
  assign _GEN_1179 = _T_599 ? buf_13_reserved : _GEN_1162; // @[ROB.scala 94:29]
  assign _GEN_1180 = _T_586 | _GEN_1179; // @[ROB.scala 92:32]
  assign _T_600 = io_graduate_0_bits_addr == 4'he; // @[ROB.scala 68:36]
  assign _T_601 = io_graduate_0_valid & _T_600; // @[ROB.scala 68:20]
  assign _T_602_valid = _T_601 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_602_bits_addr = _T_601 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_605 = _T_8_bits_addr <= 4'he; // @[ROB.scala 71:61]
  assign _T_606 = _T_16 & _T_605; // @[ROB.scala 71:41]
  assign _T_607 = 4'he < unreserved; // @[ROB.scala 71:75]
  assign _T_608 = _T_606 & _T_607; // @[ROB.scala 71:68]
  assign _T_612 = _T_607 | _T_605; // @[ROB.scala 72:61]
  assign _T_613 = _T_21 & _T_612; // @[ROB.scala 72:40]
  assign _T_614 = _T_608 | _T_613; // @[ROB.scala 71:89]
  assign _T_615 = mispredicted & _T_614; // @[ROB.scala 70:56]
  assign _T_618 = unreserved <= 4'he; // @[ROB.scala 75:55]
  assign _T_619 = 4'he < next_unreserved; // @[ROB.scala 75:69]
  assign _T_620 = _T_618 & _T_619; // @[ROB.scala 75:62]
  assign _T_621 = _T_29 & _T_620; // @[ROB.scala 75:40]
  assign _T_625 = _T_619 | _T_618; // @[ROB.scala 76:65]
  assign _T_626 = _T_34 & _T_625; // @[ROB.scala 76:39]
  assign _T_627 = _T_621 | _T_626; // @[ROB.scala 75:89]
  assign _T_628 = _T_28 & _T_627; // @[ROB.scala 74:39]
  assign _T_630 = uncommited <= 4'he; // @[ROB.scala 79:55]
  assign _T_631 = 4'he < next_uncommited; // @[ROB.scala 79:69]
  assign _T_632 = _T_630 & _T_631; // @[ROB.scala 79:62]
  assign _T_633 = _T_41 & _T_632; // @[ROB.scala 79:40]
  assign _T_637 = _T_631 | _T_630; // @[ROB.scala 80:66]
  assign _T_638 = _T_46 & _T_637; // @[ROB.scala 80:40]
  assign _T_639 = _T_633 | _T_638; // @[ROB.scala 79:89]
  assign _T_640 = _T_602_bits_addr == 4'he; // @[ROB.scala 82:60]
  assign _T_641 = _T_602_valid & _T_640; // @[ROB.scala 82:38]
  assign _GEN_1212 = _T_639 ? 1'h0 : buf_14_reserved; // @[ROB.scala 98:31]
  assign _GEN_1213 = _T_639 ? 1'h0 : buf_14_committable; // @[ROB.scala 98:31]
  assign _GEN_1214 = _T_641 | _GEN_1213; // @[ROB.scala 94:29]
  assign _GEN_1229 = _T_641 ? buf_14_reserved : _GEN_1212; // @[ROB.scala 94:29]
  assign _GEN_1230 = _T_628 | _GEN_1229; // @[ROB.scala 92:32]
  assign _T_642 = io_graduate_0_bits_addr == 4'hf; // @[ROB.scala 68:36]
  assign _T_643 = io_graduate_0_valid & _T_642; // @[ROB.scala 68:20]
  assign _T_644_valid = _T_643 ? io_graduate_0_valid : io_graduate_1_valid; // @[ROB.scala 68:10]
  assign _T_644_bits_addr = _T_643 ? io_graduate_0_bits_addr : io_graduate_1_bits_addr; // @[ROB.scala 68:10]
  assign _T_657 = mispredicted & _T_21; // @[ROB.scala 70:56]
  assign _T_670 = _T_28 & _T_34; // @[ROB.scala 74:39]
  assign _T_682 = _T_644_bits_addr == 4'hf; // @[ROB.scala 82:60]
  assign _T_683 = _T_644_valid & _T_682; // @[ROB.scala 82:38]
  assign _GEN_1262 = _T_46 ? 1'h0 : buf_15_reserved; // @[ROB.scala 98:31]
  assign _GEN_1263 = _T_46 ? 1'h0 : buf_15_committable; // @[ROB.scala 98:31]
  assign _GEN_1264 = _T_683 | _GEN_1263; // @[ROB.scala 94:29]
  assign _GEN_1279 = _T_683 ? buf_15_reserved : _GEN_1262; // @[ROB.scala 94:29]
  assign _GEN_1280 = _T_670 | _GEN_1279; // @[ROB.scala 92:32]
  assign _T_686 = 1'h0 < commitable_0; // @[ROB.scala 106:15]
  assign _GEN_1570 = _T_686 ? {{4'd0}, _GEN_240} : 20'ha00af; // @[ROB.scala 106:33]
  assign _T_689 = {{1'd0}, unreserved}; // @[ROB.scala 118:46]
  assign _T_691 = $unsigned(reset); // @[ROB.scala 121:9]
  assign _T_692 = _T_691 == 1'h0; // @[ROB.scala 121:9]
  assign io_commit_0_rd_addr = _T_686 ? _GEN_244 : 3'h0; // @[ROB.scala 108:28 ROB.scala 112:28]
  assign io_commit_0_rf_w = _T_686 & _GEN_249; // @[ROB.scala 107:25 ROB.scala 111:25]
  assign io_commit_0_data = _GEN_1570[15:0]; // @[ROB.scala 109:25 ROB.scala 113:25]
  assign io_unreserved_head_0_valid = unreserved_add_used_valid & _T_28; // @[ROB.scala 117:33]
  assign io_unreserved_head_0_bits = _T_689[3:0]; // @[ROB.scala 118:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_data = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  buf_0_inst_info_rd_addr = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  buf_0_inst_info_ctrl_rf_w = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  buf_0_reserved = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  buf_0_committable = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  buf_1_data = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  buf_1_inst_info_rd_addr = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  buf_1_inst_info_ctrl_rf_w = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  buf_1_reserved = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  buf_1_committable = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  buf_2_data = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  buf_2_inst_info_rd_addr = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  buf_2_inst_info_ctrl_rf_w = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  buf_2_reserved = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  buf_2_committable = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  buf_3_data = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  buf_3_inst_info_rd_addr = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  buf_3_inst_info_ctrl_rf_w = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  buf_3_reserved = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  buf_3_committable = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  buf_4_data = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  buf_4_inst_info_rd_addr = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  buf_4_inst_info_ctrl_rf_w = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  buf_4_reserved = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  buf_4_committable = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  buf_5_data = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  buf_5_inst_info_rd_addr = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  buf_5_inst_info_ctrl_rf_w = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  buf_5_reserved = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  buf_5_committable = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  buf_6_data = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  buf_6_inst_info_rd_addr = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  buf_6_inst_info_ctrl_rf_w = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  buf_6_reserved = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  buf_6_committable = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  buf_7_data = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  buf_7_inst_info_rd_addr = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  buf_7_inst_info_ctrl_rf_w = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  buf_7_reserved = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  buf_7_committable = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  buf_8_data = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  buf_8_inst_info_rd_addr = _RAND_41[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  buf_8_inst_info_ctrl_rf_w = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  buf_8_reserved = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  buf_8_committable = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  buf_9_data = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  buf_9_inst_info_rd_addr = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  buf_9_inst_info_ctrl_rf_w = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  buf_9_reserved = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  buf_9_committable = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  buf_10_data = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  buf_10_inst_info_rd_addr = _RAND_51[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  buf_10_inst_info_ctrl_rf_w = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  buf_10_reserved = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  buf_10_committable = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  buf_11_data = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  buf_11_inst_info_rd_addr = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  buf_11_inst_info_ctrl_rf_w = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  buf_11_reserved = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  buf_11_committable = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  buf_12_data = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  buf_12_inst_info_rd_addr = _RAND_61[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  buf_12_inst_info_ctrl_rf_w = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  buf_12_reserved = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  buf_12_committable = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  buf_13_data = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  buf_13_inst_info_rd_addr = _RAND_66[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  buf_13_inst_info_ctrl_rf_w = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  buf_13_reserved = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  buf_13_committable = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  buf_14_data = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  buf_14_inst_info_rd_addr = _RAND_71[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  buf_14_inst_info_ctrl_rf_w = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  buf_14_reserved = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  buf_14_committable = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  buf_15_data = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  buf_15_inst_info_rd_addr = _RAND_76[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  buf_15_inst_info_ctrl_rf_w = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  buf_15_reserved = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  buf_15_committable = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  uncommited = _RAND_80[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  unreserved = _RAND_81[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      buf_0_data <= 16'h0;
    end else if (!(_T_27)) begin
      if (!(_T_40)) begin
        if (_T_53) begin
          if (_T_13) begin
            buf_0_data <= io_graduate_0_bits_data;
          end else begin
            buf_0_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_0_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_27)) begin
      if (!(_T_40)) begin
        if (_T_53) begin
          if (_T_13) begin
            buf_0_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_0_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_0_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_27)) begin
      if (!(_T_40)) begin
        if (_T_53) begin
          if (_T_13) begin
            buf_0_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_0_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_0_reserved <= 1'h0;
    end else if (_T_27) begin
      buf_0_reserved <= 1'h0;
    end else begin
      buf_0_reserved <= _GEN_530;
    end
    if (reset) begin
      buf_0_committable <= 1'h0;
    end else if (_T_27) begin
      buf_0_committable <= 1'h0;
    end else if (!(_T_40)) begin
      buf_0_committable <= _GEN_514;
    end
    if (reset) begin
      buf_1_data <= 16'h0;
    end else if (!(_T_69)) begin
      if (!(_T_82)) begin
        if (_T_95) begin
          if (_T_55) begin
            buf_1_data <= io_graduate_0_bits_data;
          end else begin
            buf_1_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_1_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_69)) begin
      if (!(_T_82)) begin
        if (_T_95) begin
          if (_T_55) begin
            buf_1_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_1_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_1_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_69)) begin
      if (!(_T_82)) begin
        if (_T_95) begin
          if (_T_55) begin
            buf_1_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_1_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_1_reserved <= 1'h0;
    end else if (_T_69) begin
      buf_1_reserved <= 1'h0;
    end else begin
      buf_1_reserved <= _GEN_580;
    end
    if (reset) begin
      buf_1_committable <= 1'h0;
    end else if (_T_69) begin
      buf_1_committable <= 1'h0;
    end else if (!(_T_82)) begin
      buf_1_committable <= _GEN_564;
    end
    if (reset) begin
      buf_2_data <= 16'h0;
    end else if (!(_T_111)) begin
      if (!(_T_124)) begin
        if (_T_137) begin
          if (_T_97) begin
            buf_2_data <= io_graduate_0_bits_data;
          end else begin
            buf_2_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_2_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_111)) begin
      if (!(_T_124)) begin
        if (_T_137) begin
          if (_T_97) begin
            buf_2_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_2_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_2_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_111)) begin
      if (!(_T_124)) begin
        if (_T_137) begin
          if (_T_97) begin
            buf_2_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_2_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_2_reserved <= 1'h0;
    end else if (_T_111) begin
      buf_2_reserved <= 1'h0;
    end else begin
      buf_2_reserved <= _GEN_630;
    end
    if (reset) begin
      buf_2_committable <= 1'h0;
    end else if (_T_111) begin
      buf_2_committable <= 1'h0;
    end else if (!(_T_124)) begin
      buf_2_committable <= _GEN_614;
    end
    if (reset) begin
      buf_3_data <= 16'h0;
    end else if (!(_T_153)) begin
      if (!(_T_166)) begin
        if (_T_179) begin
          if (_T_139) begin
            buf_3_data <= io_graduate_0_bits_data;
          end else begin
            buf_3_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_3_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_153)) begin
      if (!(_T_166)) begin
        if (_T_179) begin
          if (_T_139) begin
            buf_3_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_3_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_3_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_153)) begin
      if (!(_T_166)) begin
        if (_T_179) begin
          if (_T_139) begin
            buf_3_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_3_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_3_reserved <= 1'h0;
    end else if (_T_153) begin
      buf_3_reserved <= 1'h0;
    end else begin
      buf_3_reserved <= _GEN_680;
    end
    if (reset) begin
      buf_3_committable <= 1'h0;
    end else if (_T_153) begin
      buf_3_committable <= 1'h0;
    end else if (!(_T_166)) begin
      buf_3_committable <= _GEN_664;
    end
    if (reset) begin
      buf_4_data <= 16'h0;
    end else if (!(_T_195)) begin
      if (!(_T_208)) begin
        if (_T_221) begin
          if (_T_181) begin
            buf_4_data <= io_graduate_0_bits_data;
          end else begin
            buf_4_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_4_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_195)) begin
      if (!(_T_208)) begin
        if (_T_221) begin
          if (_T_181) begin
            buf_4_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_4_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_4_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_195)) begin
      if (!(_T_208)) begin
        if (_T_221) begin
          if (_T_181) begin
            buf_4_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_4_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_4_reserved <= 1'h0;
    end else if (_T_195) begin
      buf_4_reserved <= 1'h0;
    end else begin
      buf_4_reserved <= _GEN_730;
    end
    if (reset) begin
      buf_4_committable <= 1'h0;
    end else if (_T_195) begin
      buf_4_committable <= 1'h0;
    end else if (!(_T_208)) begin
      buf_4_committable <= _GEN_714;
    end
    if (reset) begin
      buf_5_data <= 16'h0;
    end else if (!(_T_237)) begin
      if (!(_T_250)) begin
        if (_T_263) begin
          if (_T_223) begin
            buf_5_data <= io_graduate_0_bits_data;
          end else begin
            buf_5_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_5_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_237)) begin
      if (!(_T_250)) begin
        if (_T_263) begin
          if (_T_223) begin
            buf_5_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_5_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_5_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_237)) begin
      if (!(_T_250)) begin
        if (_T_263) begin
          if (_T_223) begin
            buf_5_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_5_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_5_reserved <= 1'h0;
    end else if (_T_237) begin
      buf_5_reserved <= 1'h0;
    end else begin
      buf_5_reserved <= _GEN_780;
    end
    if (reset) begin
      buf_5_committable <= 1'h0;
    end else if (_T_237) begin
      buf_5_committable <= 1'h0;
    end else if (!(_T_250)) begin
      buf_5_committable <= _GEN_764;
    end
    if (reset) begin
      buf_6_data <= 16'h0;
    end else if (!(_T_279)) begin
      if (!(_T_292)) begin
        if (_T_305) begin
          if (_T_265) begin
            buf_6_data <= io_graduate_0_bits_data;
          end else begin
            buf_6_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_6_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_279)) begin
      if (!(_T_292)) begin
        if (_T_305) begin
          if (_T_265) begin
            buf_6_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_6_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_6_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_279)) begin
      if (!(_T_292)) begin
        if (_T_305) begin
          if (_T_265) begin
            buf_6_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_6_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_6_reserved <= 1'h0;
    end else if (_T_279) begin
      buf_6_reserved <= 1'h0;
    end else begin
      buf_6_reserved <= _GEN_830;
    end
    if (reset) begin
      buf_6_committable <= 1'h0;
    end else if (_T_279) begin
      buf_6_committable <= 1'h0;
    end else if (!(_T_292)) begin
      buf_6_committable <= _GEN_814;
    end
    if (reset) begin
      buf_7_data <= 16'h0;
    end else if (!(_T_321)) begin
      if (!(_T_334)) begin
        if (_T_347) begin
          if (_T_307) begin
            buf_7_data <= io_graduate_0_bits_data;
          end else begin
            buf_7_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_7_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_321)) begin
      if (!(_T_334)) begin
        if (_T_347) begin
          if (_T_307) begin
            buf_7_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_7_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_7_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_321)) begin
      if (!(_T_334)) begin
        if (_T_347) begin
          if (_T_307) begin
            buf_7_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_7_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_7_reserved <= 1'h0;
    end else if (_T_321) begin
      buf_7_reserved <= 1'h0;
    end else begin
      buf_7_reserved <= _GEN_880;
    end
    if (reset) begin
      buf_7_committable <= 1'h0;
    end else if (_T_321) begin
      buf_7_committable <= 1'h0;
    end else if (!(_T_334)) begin
      buf_7_committable <= _GEN_864;
    end
    if (reset) begin
      buf_8_data <= 16'h0;
    end else if (!(_T_363)) begin
      if (!(_T_376)) begin
        if (_T_389) begin
          if (_T_349) begin
            buf_8_data <= io_graduate_0_bits_data;
          end else begin
            buf_8_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_8_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_363)) begin
      if (!(_T_376)) begin
        if (_T_389) begin
          if (_T_349) begin
            buf_8_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_8_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_8_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_363)) begin
      if (!(_T_376)) begin
        if (_T_389) begin
          if (_T_349) begin
            buf_8_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_8_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_8_reserved <= 1'h0;
    end else if (_T_363) begin
      buf_8_reserved <= 1'h0;
    end else begin
      buf_8_reserved <= _GEN_930;
    end
    if (reset) begin
      buf_8_committable <= 1'h0;
    end else if (_T_363) begin
      buf_8_committable <= 1'h0;
    end else if (!(_T_376)) begin
      buf_8_committable <= _GEN_914;
    end
    if (reset) begin
      buf_9_data <= 16'h0;
    end else if (!(_T_405)) begin
      if (!(_T_418)) begin
        if (_T_431) begin
          if (_T_391) begin
            buf_9_data <= io_graduate_0_bits_data;
          end else begin
            buf_9_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_9_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_405)) begin
      if (!(_T_418)) begin
        if (_T_431) begin
          if (_T_391) begin
            buf_9_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_9_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_9_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_405)) begin
      if (!(_T_418)) begin
        if (_T_431) begin
          if (_T_391) begin
            buf_9_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_9_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_9_reserved <= 1'h0;
    end else if (_T_405) begin
      buf_9_reserved <= 1'h0;
    end else begin
      buf_9_reserved <= _GEN_980;
    end
    if (reset) begin
      buf_9_committable <= 1'h0;
    end else if (_T_405) begin
      buf_9_committable <= 1'h0;
    end else if (!(_T_418)) begin
      buf_9_committable <= _GEN_964;
    end
    if (reset) begin
      buf_10_data <= 16'h0;
    end else if (!(_T_447)) begin
      if (!(_T_460)) begin
        if (_T_473) begin
          if (_T_433) begin
            buf_10_data <= io_graduate_0_bits_data;
          end else begin
            buf_10_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_10_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_447)) begin
      if (!(_T_460)) begin
        if (_T_473) begin
          if (_T_433) begin
            buf_10_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_10_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_10_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_447)) begin
      if (!(_T_460)) begin
        if (_T_473) begin
          if (_T_433) begin
            buf_10_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_10_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_10_reserved <= 1'h0;
    end else if (_T_447) begin
      buf_10_reserved <= 1'h0;
    end else begin
      buf_10_reserved <= _GEN_1030;
    end
    if (reset) begin
      buf_10_committable <= 1'h0;
    end else if (_T_447) begin
      buf_10_committable <= 1'h0;
    end else if (!(_T_460)) begin
      buf_10_committable <= _GEN_1014;
    end
    if (reset) begin
      buf_11_data <= 16'h0;
    end else if (!(_T_489)) begin
      if (!(_T_502)) begin
        if (_T_515) begin
          if (_T_475) begin
            buf_11_data <= io_graduate_0_bits_data;
          end else begin
            buf_11_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_11_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_489)) begin
      if (!(_T_502)) begin
        if (_T_515) begin
          if (_T_475) begin
            buf_11_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_11_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_11_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_489)) begin
      if (!(_T_502)) begin
        if (_T_515) begin
          if (_T_475) begin
            buf_11_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_11_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_11_reserved <= 1'h0;
    end else if (_T_489) begin
      buf_11_reserved <= 1'h0;
    end else begin
      buf_11_reserved <= _GEN_1080;
    end
    if (reset) begin
      buf_11_committable <= 1'h0;
    end else if (_T_489) begin
      buf_11_committable <= 1'h0;
    end else if (!(_T_502)) begin
      buf_11_committable <= _GEN_1064;
    end
    if (reset) begin
      buf_12_data <= 16'h0;
    end else if (!(_T_531)) begin
      if (!(_T_544)) begin
        if (_T_557) begin
          if (_T_517) begin
            buf_12_data <= io_graduate_0_bits_data;
          end else begin
            buf_12_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_12_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_531)) begin
      if (!(_T_544)) begin
        if (_T_557) begin
          if (_T_517) begin
            buf_12_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_12_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_12_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_531)) begin
      if (!(_T_544)) begin
        if (_T_557) begin
          if (_T_517) begin
            buf_12_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_12_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_12_reserved <= 1'h0;
    end else if (_T_531) begin
      buf_12_reserved <= 1'h0;
    end else begin
      buf_12_reserved <= _GEN_1130;
    end
    if (reset) begin
      buf_12_committable <= 1'h0;
    end else if (_T_531) begin
      buf_12_committable <= 1'h0;
    end else if (!(_T_544)) begin
      buf_12_committable <= _GEN_1114;
    end
    if (reset) begin
      buf_13_data <= 16'h0;
    end else if (!(_T_573)) begin
      if (!(_T_586)) begin
        if (_T_599) begin
          if (_T_559) begin
            buf_13_data <= io_graduate_0_bits_data;
          end else begin
            buf_13_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_13_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_573)) begin
      if (!(_T_586)) begin
        if (_T_599) begin
          if (_T_559) begin
            buf_13_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_13_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_13_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_573)) begin
      if (!(_T_586)) begin
        if (_T_599) begin
          if (_T_559) begin
            buf_13_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_13_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_13_reserved <= 1'h0;
    end else if (_T_573) begin
      buf_13_reserved <= 1'h0;
    end else begin
      buf_13_reserved <= _GEN_1180;
    end
    if (reset) begin
      buf_13_committable <= 1'h0;
    end else if (_T_573) begin
      buf_13_committable <= 1'h0;
    end else if (!(_T_586)) begin
      buf_13_committable <= _GEN_1164;
    end
    if (reset) begin
      buf_14_data <= 16'h0;
    end else if (!(_T_615)) begin
      if (!(_T_628)) begin
        if (_T_641) begin
          if (_T_601) begin
            buf_14_data <= io_graduate_0_bits_data;
          end else begin
            buf_14_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_14_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_615)) begin
      if (!(_T_628)) begin
        if (_T_641) begin
          if (_T_601) begin
            buf_14_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_14_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_14_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_615)) begin
      if (!(_T_628)) begin
        if (_T_641) begin
          if (_T_601) begin
            buf_14_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_14_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_14_reserved <= 1'h0;
    end else if (_T_615) begin
      buf_14_reserved <= 1'h0;
    end else begin
      buf_14_reserved <= _GEN_1230;
    end
    if (reset) begin
      buf_14_committable <= 1'h0;
    end else if (_T_615) begin
      buf_14_committable <= 1'h0;
    end else if (!(_T_628)) begin
      buf_14_committable <= _GEN_1214;
    end
    if (reset) begin
      buf_15_data <= 16'h0;
    end else if (!(_T_657)) begin
      if (!(_T_670)) begin
        if (_T_683) begin
          if (_T_643) begin
            buf_15_data <= io_graduate_0_bits_data;
          end else begin
            buf_15_data <= io_graduate_1_bits_data;
          end
        end
      end
    end
    if (reset) begin
      buf_15_inst_info_rd_addr <= 3'h0;
    end else if (!(_T_657)) begin
      if (!(_T_670)) begin
        if (_T_683) begin
          if (_T_643) begin
            buf_15_inst_info_rd_addr <= io_graduate_0_bits_inst_info_rd_addr;
          end else begin
            buf_15_inst_info_rd_addr <= io_graduate_1_bits_inst_info_rd_addr;
          end
        end
      end
    end
    if (reset) begin
      buf_15_inst_info_ctrl_rf_w <= 1'h0;
    end else if (!(_T_657)) begin
      if (!(_T_670)) begin
        if (_T_683) begin
          if (_T_643) begin
            buf_15_inst_info_ctrl_rf_w <= io_graduate_0_bits_inst_info_ctrl_rf_w;
          end else begin
            buf_15_inst_info_ctrl_rf_w <= io_graduate_1_bits_inst_info_ctrl_rf_w;
          end
        end
      end
    end
    if (reset) begin
      buf_15_reserved <= 1'h0;
    end else if (_T_657) begin
      buf_15_reserved <= 1'h0;
    end else begin
      buf_15_reserved <= _GEN_1280;
    end
    if (reset) begin
      buf_15_committable <= 1'h0;
    end else if (_T_657) begin
      buf_15_committable <= 1'h0;
    end else if (!(_T_670)) begin
      buf_15_committable <= _GEN_1264;
    end
    if (reset) begin
      uncommited <= 4'h0;
    end else begin
      uncommited <= next_uncommited;
    end
    if (reset) begin
      unreserved <= 4'h0;
    end else if (mispredicted) begin
      if (_T_7) begin
        unreserved <= io_graduate_0_bits_addr;
      end else begin
        unreserved <= io_graduate_1_bits_addr;
      end
    end else if (unreserved_add_used_valid) begin
      unreserved <= unreserved_add_used;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_692) begin
          $fwrite(32'h80000002,"unreserved: %d, next_unreserved: %d\n",unreserved,next_unreserved); // @[ROB.scala 121:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_692) begin
          $fwrite(32'h80000002,"uncommited: %d, next_uncommited: %d, can_commit_cnt: %d\n",uncommited,next_uncommited,commitable_0); // @[ROB.scala 122:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_692) begin
          $fwrite(32'h80000002,"mispredicted: %d, unreserved_add_used_valid: %d\n",mispredicted,unreserved_add_used_valid); // @[ROB.scala 123:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_692) begin
          $fwrite(32'h80000002,"-----------------------------------\n"); // @[ROB.scala 124:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Hart(
  input         clock,
  input         reset,
  output [15:0] io_pc,
  output [15:0] io_total_cnt,
  output [15:0] io_rf_0,
  output [15:0] io_rf_1,
  output [15:0] io_rf_2,
  output [15:0] io_rf_3,
  output [15:0] io_rf_4,
  output [15:0] io_rf_5,
  output [15:0] io_rf_6,
  output [15:0] io_rf_7
);
  wire  m_bp_clock; // @[Hart.scala 36:37]
  wire  m_bp_reset; // @[Hart.scala 36:37]
  wire [15:0] m_bp_io_pc; // @[Hart.scala 36:37]
  wire  m_bp_io_stall; // @[Hart.scala 36:37]
  wire  m_bp_io_learning_valid; // @[Hart.scala 36:37]
  wire [15:0] m_bp_io_learning_bits_pc; // @[Hart.scala 36:37]
  wire  m_bp_io_learning_bits_result; // @[Hart.scala 36:37]
  wire  m_bp_io_predict; // @[Hart.scala 36:37]
  wire  s_if_clock; // @[Hart.scala 37:24]
  wire  s_if_reset; // @[Hart.scala 37:24]
  wire  s_if_io_in_branch_mispredicted; // @[Hart.scala 37:24]
  wire  s_if_io_in_branch_graduated; // @[Hart.scala 37:24]
  wire [15:0] s_if_io_in_restoration_pc; // @[Hart.scala 37:24]
  wire  s_if_io_in_predict; // @[Hart.scala 37:24]
  wire  s_if_io_in_predict_enable; // @[Hart.scala 37:24]
  wire [15:0] s_if_io_in_predict_pc; // @[Hart.scala 37:24]
  wire  s_if_io_in_is_jump; // @[Hart.scala 37:24]
  wire [15:0] s_if_io_in_jump_pc; // @[Hart.scala 37:24]
  wire  s_if_io_in_stall; // @[Hart.scala 37:24]
  wire [15:0] s_if_io_out_pc; // @[Hart.scala 37:24]
  wire [15:0] s_if_io_out_total_cnt; // @[Hart.scala 37:24]
  wire [3:0] s_if_io_out_inst_bits_op; // @[Hart.scala 37:24]
  wire [2:0] s_if_io_out_inst_bits_rd; // @[Hart.scala 37:24]
  wire [2:0] s_if_io_out_inst_bits_rs; // @[Hart.scala 37:24]
  wire [5:0] s_if_io_out_inst_bits_disp6u; // @[Hart.scala 37:24]
  wire  s_id_clock; // @[Hart.scala 38:24]
  wire  s_id_reset; // @[Hart.scala 38:24]
  wire  s_id_io_predict; // @[Hart.scala 38:24]
  wire  s_id_io_branch_mispredicted; // @[Hart.scala 38:24]
  wire  s_id_io_branch_graduated; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_if_out_pc; // @[Hart.scala 38:24]
  wire [3:0] s_id_io_if_out_inst_bits_op; // @[Hart.scala 38:24]
  wire [2:0] s_id_io_if_out_inst_bits_rd; // @[Hart.scala 38:24]
  wire [2:0] s_id_io_if_out_inst_bits_rs; // @[Hart.scala 38:24]
  wire [5:0] s_id_io_if_out_inst_bits_disp6u; // @[Hart.scala 38:24]
  wire [2:0] s_id_io_commit_0_rd_addr; // @[Hart.scala 38:24]
  wire  s_id_io_commit_0_rf_w; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_commit_0_data; // @[Hart.scala 38:24]
  wire  s_id_io_unreserved_head_0_valid; // @[Hart.scala 38:24]
  wire [3:0] s_id_io_unreserved_head_0_bits; // @[Hart.scala 38:24]
  wire  s_id_io_used_num; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_jump_pc; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_next_pc; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_valid; // @[Hart.scala 38:24]
  wire [2:0] s_id_io_inst_info_rd_addr; // @[Hart.scala 38:24]
  wire [3:0] s_id_io_inst_info_rob_addr; // @[Hart.scala 38:24]
  wire [2:0] s_id_io_inst_info_ctrl_alu_op; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_ctrl_is_jump; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_ctrl_is_branch; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_ctrl_rf_w; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_ctrl_mem_r; // @[Hart.scala 38:24]
  wire  s_id_io_inst_info_ctrl_mem_w; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_source_0; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_source_1; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rd; // @[Hart.scala 38:24]
  wire  s_id_io_stall; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_pc; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_1; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_2; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_3; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_4; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_5; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_6; // @[Hart.scala 38:24]
  wire [15:0] s_id_io_rf4debug_7; // @[Hart.scala 38:24]
  wire  s_ex_clock; // @[Hart.scala 39:24]
  wire  s_ex_reset; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_valid; // @[Hart.scala 39:24]
  wire [2:0] s_ex_io_inst_info_rd_addr; // @[Hart.scala 39:24]
  wire [3:0] s_ex_io_inst_info_rob_addr; // @[Hart.scala 39:24]
  wire [2:0] s_ex_io_inst_info_ctrl_alu_op; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_ctrl_is_branch; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_ctrl_rf_w; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_ctrl_mem_r; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_ctrl_mem_w; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_source_0; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_source_1; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_branch_pc; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_next_pc; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_rd; // @[Hart.scala 39:24]
  wire  s_ex_io_predict; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_pc; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_alu_out; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_out_valid; // @[Hart.scala 39:24]
  wire [2:0] s_ex_io_inst_info_out_rd_addr; // @[Hart.scala 39:24]
  wire [3:0] s_ex_io_inst_info_out_rob_addr; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_out_ctrl_is_branch; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_out_ctrl_rf_w; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_out_ctrl_mem_r; // @[Hart.scala 39:24]
  wire  s_ex_io_inst_info_out_ctrl_mem_w; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_restoration_pc_out; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_rd_out; // @[Hart.scala 39:24]
  wire [15:0] s_ex_io_pc_out; // @[Hart.scala 39:24]
  wire  s_ex_io_mispredicted; // @[Hart.scala 39:24]
  wire  s_im_clock; // @[Hart.scala 40:24]
  wire  s_im_io_inst_info_valid; // @[Hart.scala 40:24]
  wire [2:0] s_im_io_inst_info_rd_addr; // @[Hart.scala 40:24]
  wire [3:0] s_im_io_inst_info_rob_addr; // @[Hart.scala 40:24]
  wire  s_im_io_inst_info_ctrl_rf_w; // @[Hart.scala 40:24]
  wire  s_im_io_inst_info_ctrl_mem_r; // @[Hart.scala 40:24]
  wire  s_im_io_inst_info_ctrl_mem_w; // @[Hart.scala 40:24]
  wire [3:0] s_im_io_rd_out; // @[Hart.scala 40:24]
  wire [3:0] s_im_io_alu_out; // @[Hart.scala 40:24]
  wire [15:0] s_im_io_mem_out; // @[Hart.scala 40:24]
  wire  m_rob_clock; // @[Hart.scala 41:26]
  wire  m_rob_reset; // @[Hart.scala 41:26]
  wire  m_rob_io_used_num; // @[Hart.scala 41:26]
  wire  m_rob_io_graduate_0_valid; // @[Hart.scala 41:26]
  wire [15:0] m_rob_io_graduate_0_bits_data; // @[Hart.scala 41:26]
  wire [2:0] m_rob_io_graduate_0_bits_inst_info_rd_addr; // @[Hart.scala 41:26]
  wire  m_rob_io_graduate_0_bits_inst_info_ctrl_rf_w; // @[Hart.scala 41:26]
  wire [3:0] m_rob_io_graduate_0_bits_addr; // @[Hart.scala 41:26]
  wire  m_rob_io_graduate_0_bits_mispredicted; // @[Hart.scala 41:26]
  wire  m_rob_io_graduate_1_valid; // @[Hart.scala 41:26]
  wire [15:0] m_rob_io_graduate_1_bits_data; // @[Hart.scala 41:26]
  wire [2:0] m_rob_io_graduate_1_bits_inst_info_rd_addr; // @[Hart.scala 41:26]
  wire  m_rob_io_graduate_1_bits_inst_info_ctrl_rf_w; // @[Hart.scala 41:26]
  wire [3:0] m_rob_io_graduate_1_bits_addr; // @[Hart.scala 41:26]
  wire [2:0] m_rob_io_commit_0_rd_addr; // @[Hart.scala 41:26]
  wire  m_rob_io_commit_0_rf_w; // @[Hart.scala 41:26]
  wire [15:0] m_rob_io_commit_0_data; // @[Hart.scala 41:26]
  wire  m_rob_io_unreserved_head_0_valid; // @[Hart.scala 41:26]
  wire [3:0] m_rob_io_unreserved_head_0_bits; // @[Hart.scala 41:26]
  BranchPredictor m_bp ( // @[Hart.scala 36:37]
    .clock(m_bp_clock),
    .reset(m_bp_reset),
    .io_pc(m_bp_io_pc),
    .io_stall(m_bp_io_stall),
    .io_learning_valid(m_bp_io_learning_valid),
    .io_learning_bits_pc(m_bp_io_learning_bits_pc),
    .io_learning_bits_result(m_bp_io_learning_bits_result),
    .io_predict(m_bp_io_predict)
  );
  IF s_if ( // @[Hart.scala 37:24]
    .clock(s_if_clock),
    .reset(s_if_reset),
    .io_in_branch_mispredicted(s_if_io_in_branch_mispredicted),
    .io_in_branch_graduated(s_if_io_in_branch_graduated),
    .io_in_restoration_pc(s_if_io_in_restoration_pc),
    .io_in_predict(s_if_io_in_predict),
    .io_in_predict_enable(s_if_io_in_predict_enable),
    .io_in_predict_pc(s_if_io_in_predict_pc),
    .io_in_is_jump(s_if_io_in_is_jump),
    .io_in_jump_pc(s_if_io_in_jump_pc),
    .io_in_stall(s_if_io_in_stall),
    .io_out_pc(s_if_io_out_pc),
    .io_out_total_cnt(s_if_io_out_total_cnt),
    .io_out_inst_bits_op(s_if_io_out_inst_bits_op),
    .io_out_inst_bits_rd(s_if_io_out_inst_bits_rd),
    .io_out_inst_bits_rs(s_if_io_out_inst_bits_rs),
    .io_out_inst_bits_disp6u(s_if_io_out_inst_bits_disp6u)
  );
  ID s_id ( // @[Hart.scala 38:24]
    .clock(s_id_clock),
    .reset(s_id_reset),
    .io_predict(s_id_io_predict),
    .io_branch_mispredicted(s_id_io_branch_mispredicted),
    .io_branch_graduated(s_id_io_branch_graduated),
    .io_if_out_pc(s_id_io_if_out_pc),
    .io_if_out_inst_bits_op(s_id_io_if_out_inst_bits_op),
    .io_if_out_inst_bits_rd(s_id_io_if_out_inst_bits_rd),
    .io_if_out_inst_bits_rs(s_id_io_if_out_inst_bits_rs),
    .io_if_out_inst_bits_disp6u(s_id_io_if_out_inst_bits_disp6u),
    .io_commit_0_rd_addr(s_id_io_commit_0_rd_addr),
    .io_commit_0_rf_w(s_id_io_commit_0_rf_w),
    .io_commit_0_data(s_id_io_commit_0_data),
    .io_unreserved_head_0_valid(s_id_io_unreserved_head_0_valid),
    .io_unreserved_head_0_bits(s_id_io_unreserved_head_0_bits),
    .io_used_num(s_id_io_used_num),
    .io_jump_pc(s_id_io_jump_pc),
    .io_next_pc(s_id_io_next_pc),
    .io_inst_info_valid(s_id_io_inst_info_valid),
    .io_inst_info_rd_addr(s_id_io_inst_info_rd_addr),
    .io_inst_info_rob_addr(s_id_io_inst_info_rob_addr),
    .io_inst_info_ctrl_alu_op(s_id_io_inst_info_ctrl_alu_op),
    .io_inst_info_ctrl_is_jump(s_id_io_inst_info_ctrl_is_jump),
    .io_inst_info_ctrl_is_branch(s_id_io_inst_info_ctrl_is_branch),
    .io_inst_info_ctrl_rf_w(s_id_io_inst_info_ctrl_rf_w),
    .io_inst_info_ctrl_mem_r(s_id_io_inst_info_ctrl_mem_r),
    .io_inst_info_ctrl_mem_w(s_id_io_inst_info_ctrl_mem_w),
    .io_source_0(s_id_io_source_0),
    .io_source_1(s_id_io_source_1),
    .io_rd(s_id_io_rd),
    .io_stall(s_id_io_stall),
    .io_pc(s_id_io_pc),
    .io_rf4debug_1(s_id_io_rf4debug_1),
    .io_rf4debug_2(s_id_io_rf4debug_2),
    .io_rf4debug_3(s_id_io_rf4debug_3),
    .io_rf4debug_4(s_id_io_rf4debug_4),
    .io_rf4debug_5(s_id_io_rf4debug_5),
    .io_rf4debug_6(s_id_io_rf4debug_6),
    .io_rf4debug_7(s_id_io_rf4debug_7)
  );
  EX s_ex ( // @[Hart.scala 39:24]
    .clock(s_ex_clock),
    .reset(s_ex_reset),
    .io_inst_info_valid(s_ex_io_inst_info_valid),
    .io_inst_info_rd_addr(s_ex_io_inst_info_rd_addr),
    .io_inst_info_rob_addr(s_ex_io_inst_info_rob_addr),
    .io_inst_info_ctrl_alu_op(s_ex_io_inst_info_ctrl_alu_op),
    .io_inst_info_ctrl_is_branch(s_ex_io_inst_info_ctrl_is_branch),
    .io_inst_info_ctrl_rf_w(s_ex_io_inst_info_ctrl_rf_w),
    .io_inst_info_ctrl_mem_r(s_ex_io_inst_info_ctrl_mem_r),
    .io_inst_info_ctrl_mem_w(s_ex_io_inst_info_ctrl_mem_w),
    .io_source_0(s_ex_io_source_0),
    .io_source_1(s_ex_io_source_1),
    .io_branch_pc(s_ex_io_branch_pc),
    .io_next_pc(s_ex_io_next_pc),
    .io_rd(s_ex_io_rd),
    .io_predict(s_ex_io_predict),
    .io_pc(s_ex_io_pc),
    .io_alu_out(s_ex_io_alu_out),
    .io_inst_info_out_valid(s_ex_io_inst_info_out_valid),
    .io_inst_info_out_rd_addr(s_ex_io_inst_info_out_rd_addr),
    .io_inst_info_out_rob_addr(s_ex_io_inst_info_out_rob_addr),
    .io_inst_info_out_ctrl_is_branch(s_ex_io_inst_info_out_ctrl_is_branch),
    .io_inst_info_out_ctrl_rf_w(s_ex_io_inst_info_out_ctrl_rf_w),
    .io_inst_info_out_ctrl_mem_r(s_ex_io_inst_info_out_ctrl_mem_r),
    .io_inst_info_out_ctrl_mem_w(s_ex_io_inst_info_out_ctrl_mem_w),
    .io_restoration_pc_out(s_ex_io_restoration_pc_out),
    .io_rd_out(s_ex_io_rd_out),
    .io_pc_out(s_ex_io_pc_out),
    .io_mispredicted(s_ex_io_mispredicted)
  );
  IM s_im ( // @[Hart.scala 40:24]
    .clock(s_im_clock),
    .io_inst_info_valid(s_im_io_inst_info_valid),
    .io_inst_info_rd_addr(s_im_io_inst_info_rd_addr),
    .io_inst_info_rob_addr(s_im_io_inst_info_rob_addr),
    .io_inst_info_ctrl_rf_w(s_im_io_inst_info_ctrl_rf_w),
    .io_inst_info_ctrl_mem_r(s_im_io_inst_info_ctrl_mem_r),
    .io_inst_info_ctrl_mem_w(s_im_io_inst_info_ctrl_mem_w),
    .io_rd_out(s_im_io_rd_out),
    .io_alu_out(s_im_io_alu_out),
    .io_mem_out(s_im_io_mem_out)
  );
  ROB m_rob ( // @[Hart.scala 41:26]
    .clock(m_rob_clock),
    .reset(m_rob_reset),
    .io_used_num(m_rob_io_used_num),
    .io_graduate_0_valid(m_rob_io_graduate_0_valid),
    .io_graduate_0_bits_data(m_rob_io_graduate_0_bits_data),
    .io_graduate_0_bits_inst_info_rd_addr(m_rob_io_graduate_0_bits_inst_info_rd_addr),
    .io_graduate_0_bits_inst_info_ctrl_rf_w(m_rob_io_graduate_0_bits_inst_info_ctrl_rf_w),
    .io_graduate_0_bits_addr(m_rob_io_graduate_0_bits_addr),
    .io_graduate_0_bits_mispredicted(m_rob_io_graduate_0_bits_mispredicted),
    .io_graduate_1_valid(m_rob_io_graduate_1_valid),
    .io_graduate_1_bits_data(m_rob_io_graduate_1_bits_data),
    .io_graduate_1_bits_inst_info_rd_addr(m_rob_io_graduate_1_bits_inst_info_rd_addr),
    .io_graduate_1_bits_inst_info_ctrl_rf_w(m_rob_io_graduate_1_bits_inst_info_ctrl_rf_w),
    .io_graduate_1_bits_addr(m_rob_io_graduate_1_bits_addr),
    .io_commit_0_rd_addr(m_rob_io_commit_0_rd_addr),
    .io_commit_0_rf_w(m_rob_io_commit_0_rf_w),
    .io_commit_0_data(m_rob_io_commit_0_data),
    .io_unreserved_head_0_valid(m_rob_io_unreserved_head_0_valid),
    .io_unreserved_head_0_bits(m_rob_io_unreserved_head_0_bits)
  );
  assign io_pc = s_if_io_out_pc; // @[Hart.scala 113:9]
  assign io_total_cnt = s_if_io_out_total_cnt; // @[Hart.scala 114:16]
  assign io_rf_0 = 16'h0; // @[Hart.scala 115:9]
  assign io_rf_1 = s_id_io_rf4debug_1; // @[Hart.scala 115:9]
  assign io_rf_2 = s_id_io_rf4debug_2; // @[Hart.scala 115:9]
  assign io_rf_3 = s_id_io_rf4debug_3; // @[Hart.scala 115:9]
  assign io_rf_4 = s_id_io_rf4debug_4; // @[Hart.scala 115:9]
  assign io_rf_5 = s_id_io_rf4debug_5; // @[Hart.scala 115:9]
  assign io_rf_6 = s_id_io_rf4debug_6; // @[Hart.scala 115:9]
  assign io_rf_7 = s_id_io_rf4debug_7; // @[Hart.scala 115:9]
  assign m_bp_clock = clock;
  assign m_bp_reset = reset;
  assign m_bp_io_pc = s_if_io_out_pc; // @[Hart.scala 61:14]
  assign m_bp_io_stall = s_id_io_stall; // @[Hart.scala 62:17]
  assign m_bp_io_learning_valid = s_ex_io_inst_info_out_ctrl_is_branch; // @[Hart.scala 63:26]
  assign m_bp_io_learning_bits_pc = s_ex_io_pc_out; // @[Hart.scala 65:28]
  assign m_bp_io_learning_bits_result = s_ex_io_alu_out[0]; // @[Hart.scala 64:32]
  assign s_if_clock = clock;
  assign s_if_reset = reset;
  assign s_if_io_in_branch_mispredicted = s_ex_io_mispredicted; // @[Hart.scala 50:34]
  assign s_if_io_in_branch_graduated = s_ex_io_inst_info_out_ctrl_is_branch; // @[Hart.scala 51:31]
  assign s_if_io_in_restoration_pc = s_ex_io_restoration_pc_out; // @[Hart.scala 52:29]
  assign s_if_io_in_predict = m_bp_io_predict; // @[Hart.scala 46:22]
  assign s_if_io_in_predict_enable = s_id_io_inst_info_ctrl_is_branch; // @[Hart.scala 47:29]
  assign s_if_io_in_predict_pc = s_id_io_jump_pc; // @[Hart.scala 48:25]
  assign s_if_io_in_is_jump = s_id_io_inst_info_ctrl_is_jump; // @[Hart.scala 54:22]
  assign s_if_io_in_jump_pc = s_id_io_jump_pc; // @[Hart.scala 55:22]
  assign s_if_io_in_stall = s_id_io_stall; // @[Hart.scala 57:20]
  assign s_id_clock = clock;
  assign s_id_reset = reset;
  assign s_id_io_predict = m_bp_io_predict; // @[Hart.scala 69:19]
  assign s_id_io_branch_mispredicted = s_ex_io_mispredicted; // @[Hart.scala 70:31]
  assign s_id_io_branch_graduated = s_ex_io_inst_info_out_ctrl_is_branch; // @[Hart.scala 71:28]
  assign s_id_io_if_out_pc = s_if_io_out_pc; // @[Hart.scala 72:18]
  assign s_id_io_if_out_inst_bits_op = s_if_io_out_inst_bits_op; // @[Hart.scala 72:18]
  assign s_id_io_if_out_inst_bits_rd = s_if_io_out_inst_bits_rd; // @[Hart.scala 72:18]
  assign s_id_io_if_out_inst_bits_rs = s_if_io_out_inst_bits_rs; // @[Hart.scala 72:18]
  assign s_id_io_if_out_inst_bits_disp6u = s_if_io_out_inst_bits_disp6u; // @[Hart.scala 72:18]
  assign s_id_io_commit_0_rd_addr = m_rob_io_commit_0_rd_addr; // @[Hart.scala 77:21]
  assign s_id_io_commit_0_rf_w = m_rob_io_commit_0_rf_w; // @[Hart.scala 77:21]
  assign s_id_io_commit_0_data = m_rob_io_commit_0_data; // @[Hart.scala 77:21]
  assign s_id_io_unreserved_head_0_valid = m_rob_io_unreserved_head_0_valid; // @[Hart.scala 79:27]
  assign s_id_io_unreserved_head_0_bits = m_rob_io_unreserved_head_0_bits; // @[Hart.scala 79:27]
  assign s_ex_clock = clock;
  assign s_ex_reset = reset;
  assign s_ex_io_inst_info_valid = s_id_io_inst_info_valid; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_rd_addr = s_id_io_inst_info_rd_addr; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_rob_addr = s_id_io_inst_info_rob_addr; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_ctrl_alu_op = s_id_io_inst_info_ctrl_alu_op; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_ctrl_is_branch = s_id_io_inst_info_ctrl_is_branch; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_ctrl_rf_w = s_id_io_inst_info_ctrl_rf_w; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_ctrl_mem_r = s_id_io_inst_info_ctrl_mem_r; // @[Hart.scala 84:21]
  assign s_ex_io_inst_info_ctrl_mem_w = s_id_io_inst_info_ctrl_mem_w; // @[Hart.scala 84:21]
  assign s_ex_io_source_0 = s_id_io_source_0; // @[Hart.scala 85:18]
  assign s_ex_io_source_1 = s_id_io_source_1; // @[Hart.scala 85:18]
  assign s_ex_io_branch_pc = s_id_io_jump_pc; // @[Hart.scala 88:21]
  assign s_ex_io_next_pc = s_id_io_next_pc; // @[Hart.scala 87:19]
  assign s_ex_io_rd = s_id_io_rd; // @[Hart.scala 86:14]
  assign s_ex_io_predict = m_bp_io_predict; // @[Hart.scala 83:19]
  assign s_ex_io_pc = s_id_io_pc; // @[Hart.scala 89:14]
  assign s_im_clock = clock;
  assign s_im_io_inst_info_valid = s_ex_io_inst_info_out_valid; // @[Hart.scala 93:21]
  assign s_im_io_inst_info_rd_addr = s_ex_io_inst_info_out_rd_addr; // @[Hart.scala 93:21]
  assign s_im_io_inst_info_rob_addr = s_ex_io_inst_info_out_rob_addr; // @[Hart.scala 93:21]
  assign s_im_io_inst_info_ctrl_rf_w = s_ex_io_inst_info_out_ctrl_rf_w; // @[Hart.scala 93:21]
  assign s_im_io_inst_info_ctrl_mem_r = s_ex_io_inst_info_out_ctrl_mem_r; // @[Hart.scala 93:21]
  assign s_im_io_inst_info_ctrl_mem_w = s_ex_io_inst_info_out_ctrl_mem_w; // @[Hart.scala 93:21]
  assign s_im_io_rd_out = s_ex_io_rd_out[3:0]; // @[Hart.scala 95:18]
  assign s_im_io_alu_out = s_ex_io_alu_out[3:0]; // @[Hart.scala 94:19]
  assign m_rob_clock = clock;
  assign m_rob_reset = reset;
  assign m_rob_io_used_num = s_id_io_used_num; // @[Hart.scala 99:21]
  assign m_rob_io_graduate_0_valid = s_ex_io_inst_info_out_valid; // @[Hart.scala 100:30]
  assign m_rob_io_graduate_0_bits_data = s_ex_io_alu_out; // @[Hart.scala 104:34]
  assign m_rob_io_graduate_0_bits_inst_info_rd_addr = s_ex_io_inst_info_out_rd_addr; // @[Hart.scala 103:39]
  assign m_rob_io_graduate_0_bits_inst_info_ctrl_rf_w = s_ex_io_inst_info_out_ctrl_rf_w; // @[Hart.scala 103:39]
  assign m_rob_io_graduate_0_bits_addr = s_ex_io_inst_info_out_rob_addr; // @[Hart.scala 101:34]
  assign m_rob_io_graduate_0_bits_mispredicted = s_ex_io_mispredicted; // @[Hart.scala 102:42]
  assign m_rob_io_graduate_1_valid = s_im_io_inst_info_valid; // @[Hart.scala 105:30]
  assign m_rob_io_graduate_1_bits_data = s_im_io_mem_out; // @[Hart.scala 109:34]
  assign m_rob_io_graduate_1_bits_inst_info_rd_addr = s_im_io_inst_info_rd_addr; // @[Hart.scala 108:39]
  assign m_rob_io_graduate_1_bits_inst_info_ctrl_rf_w = s_im_io_inst_info_ctrl_rf_w; // @[Hart.scala 108:39]
  assign m_rob_io_graduate_1_bits_addr = s_im_io_inst_info_rob_addr; // @[Hart.scala 106:34]
endmodule
